UZdnsLrj3r/HVFHPTJuK8pSMjQQXxQqlTEauDMxtQWrvlyxTCNAkMJKs/lzjBw740Cf84QsCemTP
uAYNj11KnuXF1SxW1MY2tNkOhTj2Qh6BaBLOHHNp0S8HJNW0XJykOKjHyLL98V3VpuKsHPLkKjFQ
8YqL/eybWtsTAaiyEqc1mVdywSDKyi6TNQa+RH9d6RJOH4T/nfRS4zE0c/vAXXNqb/2SEn/URkNS
M7QuJ96iyFXhtkNaAtNdI0mJT6S0OK4NZCktmITCsoyBbrSk0ZReV87Y8qMKmJhnnJ7RrX0pkALB
/0JascDxhZy/HrUcA5C4CT/2+GSC3Hjvdjt2EpSwWf+OedUaggABhX6meMSiKz7dtrByYh5Ucrv8
5kDBpAjMPWwPbd4WesnhLjQ8bQZFqajSoRqEimAM74ZuG3ov/CpAZyZcubcf9R6GZRkSb+IDqMak
k66IvK335xu3reQuNrVLrXRTTxpsovKYuGqYrizbYrg+bxCS1m2v8EEXh+/MUrRSUgTuFeHnaR32
kQDwCJlzBbdeFMugPdyS3012SxOe4Op3jW3Wdz2rnfAcvQPBXXWXffLKUunFnpW4sdFtmHqF1+Rs
can9baZxl3r9YR4dhAETZIIpfCiS4NGSILdtK0DJR1zZ92OHgnJsJaHc0/pCzs8Z5GqdO8Qm+a0/
HwGK3q7bS5yDmOC+fCRc26j4PPa9/L8tzwRhkhl+pOiYAmNjI0SuB8N4zb3kVURMlnTQfeIxWYRA
kkzCy4GmZtcf3xrX1AqTUsee2AE0jJJr6XLIJvGK26t/GbyTmZ7avo9uzSQk4S6aBQINze5fRi8r
IiDipnULdNP2YnV/1x5vP2L5nbMNsrHYIjtIIsOQR89o4bOYV55doE/8mrRNgwKhYh1sa/gjuJxJ
bSJrN5kM+mVvQLPr0QYG8JnCmU3iOSp+cEZmAAX3Hn/V9Vh2Qo+OdN4UDTEaB+Q3c14pszeqh93Y
RleDaWb73/TMcyaFUeSY/RFIBMVecWllO20ukPhuXb4FtZM222WpBB3m4/ZtXHeuTOhneulr8C7b
pNXLj7MdWMyh/fCoq6sbZaz2InPd5/yBLWXWjMe47FTnh/LHT5nwOjQR6ktSyS/k0qTonsR72vzj
ztyhvEUm9bjHEhJetfaJ/bPlLZhhgoMqYjE55Pdn5fxH731KUQ5jEGo99ePEMm60KlJDQ+/c4gSE
bqz9j0wtHU7J7orB1irq8IAyNVvUIXOTxVsQnDpXCt6VNsqKAPK6phW4KRfEzrZp3V2rhgoiyBRo
YI2BNNjwH0mOyyatGUD1Igf2ZQX/Fc1JBfSL+DcLjkDBfTLKX0Vp8+wCyHc5t6IyXw4E2dOe4VZK
w7lc+m+b5fXSfFLxCb8DxusQDpUWRCHk+ojDrMvrcAnP0bDVpwYMTYZ/qDQYzfDEa9bPHgN9WXbN
AqbTskXxrOp/HxqaAbYIkhS12QD3///DPvgcj4D/AVljDN8zFOT1B4Du3iTJpxc5cyyIvcLrYKmW
ftr1+IX2sMx3eBc9cyZ+0/6KeVR2xcbcnDLpBQKW5r0M617w8cOoMNOB/YD1wuSWw2oCC6KUS9hL
Befjio9KWxp0yEk9j3yn8sKY64AsIIgWCKkuuKy9aMiJnEQ9UYadXn5fY5h4+B0QUMNOKLVvECuG
5c8hqkJ1Y3Jv2+3kRr0+GVQtdIkBHImPpNpLFbkrjOE2wbVT7FMSJ4st3Sm5PpSEzGSCIAfbnMcz
CnZXL/7jT+NDqErDlfeYPH8iKBWDd1k2NO9b4ucfyN8Ksr5YW7LmDCzvKZjE/PH/IEgKNtpKrXVa
DoVCzT7/+AltpgcUIFirasDdQ0IfwNWtISwHWCP+kKeI4ZEg9+zIinF2xTAMfNd0uls5yY7VARhT
p3xfUEd+BBCojNNKfSu9Jop+1OHtAUqJz5TSIFZHxBAfpKsaqf9HHr1dHW7Z+cTdgdnv7aLv2ZBG
+HYHDuZqQJXsmGpOcsdOsoS8+lsEcEu4h7WZv2RKqSlkty/6PPF+WCf8xO9roJltqXo9Edb9qaj5
P0WJZCLUX7vsPmr4uedxfQMEdBqS0WlW0V/AjLlPDn6abIOZphHXUMM46RvTEFXwJQ+5S5rZJb0t
RhV3HKJgtD76QPbkNy+KOQgs2AaJbz0mdSFWFCYJLqm6T7lRLslfCfGgU3UXEbj/9TYQBBiIEYNu
tzNmTbivNlQM8OjkuwLlbsFeQq99nZlBnq46HPNHUHGXs/3eY4UxPnFC233nMaSjDe5yDJmt7KNs
MgFBJG0WvfsioktuXjYEt8lzIGtyVsPxBEpvDioBhbF3bPX8bKO9RrGiaiVljcOv3qybENdObkhZ
ch1V1YcrkM3BjNfSTc2X2DLQmEc/xe3T5iMw02zHf+tWMo0wc0WzBg3vP/N58/6hJfhwbyJSMYJD
WVpidPKqOVfIjIiMS1PPgHQLPg7GxNdOjMnVnv+Evx3m8I2KldA4EcQg3WX5xcok7yAcWhvckOud
iPDmmmrPtSb+dmJVLahsGNOCR1CwAgwNmRi/NoLUworafyEhKK1eC8jXGVwOkIyQ4J+ZnnsjbFJ6
oheAkLQXAbK7ixbwAjFEa18qNcCZ9lzK96gDTxTa7Ef3pPQOja9CjXn67suBZCTqkoKA0zWhOchz
O6u7Y0Dhy61U9tYiibBrDCuCHzAelw7pD03qbjwR9pAtsai09iI7+iTP0ZP2BQqcOlK63zi/qv+A
Q/9G+9Lby9GytObxFSrdFY76XIjrLPeo/wwDeSXTkxjBKjFzaVM9ZezFln+FzmTx1OzlmNnlJKXD
oE6CFJQjiSp7UDGWjxdhtsvJJvbLUh6lLQP1W+NjpMvUcdgShgHtSMHLqnzJD54CsBP+qp49PGUE
RXn25MdF9On6I/mMkWzTD418gCW3ywiMwoXKD/rh5rckxiujJxKQCAqQJ/g0iTp3ZRX5zmjE0lYD
ke29Z5YhnVIxaIXiQ6WnVZxgmSNvTZ2ODQNImWE0PyOZwN+McuAqE2T3cvNpFUvCuHxnsp/mWCGh
KTLdtc3OCnHNPRl7yiApd6YCVKM1G2RlzNo3auO5mm14ZXBZBJ43Q7cJySKXqcbcYRiw1VgiVwA4
VUYOtkbF2yTQDwsf9sl5uiS8s44bWlxCkXCEllC5f/O74n/+Hkmt4RBg0IY2EzuGP0vbcGudRUpa
yvYjylvqd4JQQFM6VjsMeR1T3pS7M65+DBEYu//rslLmTsU2vuf3aEJlDZL5jDl+CaaZQS3t9OHk
h4lUE2o9ZQvY4RsUOF4dOnF6gTeP51iBDwE4qmX1kqp6nafAn2Apn6bDQNTkqfxsD54y1NB97Mmo
uPIAccqylDbcpH245cbngNf8J0XnCLux19wrm8LPy85ti8pIwTkrrUeCqB2GbgnuRZ55phhWb7tu
yFCegtXjdaTDzzUjbtPGDzCdtLpRlLO1x8y1RTnW8DcKK3E5IQnKDc+MN814bw/qI2TssTFImtSr
cfgJ01qnLZIsEYJ2A49w54zSfsw8B3mG9zW62TIRJmlch0HsGm6gvbF5dyygH+aSE+bGzqktmybs
LVOnN8Hh5Xljq7xIBLadV7KTJduU2BpqlCZdXdM70aMje8GoDQd10x6J05ytcep0aPmD6PrB3haB
cpmJirTPIEPrQWbS4ZE3d3a48FeletfNDNXSY/LaUMUeYOViNBKsS20YHEd06bqQU7v9ABDe0dex
G9G91YjYuDwxje4MlSudi9TjUW+ug1GdIOAnsUmzAX8T6atOrUjhqM7TB4OS79CNo0nBWCKxO/7G
ClNlvn3yFuxmfq8lY2wxYo6F4AiJkZPXXm9CWBc60h6LCmtoxsvJOSDTfmSCOY9aykC+t0IgMKJl
TXhLE7FVAqt5GDym8mh/imjTQKeYN2PRktGoL5wrP2cCWcuQP6Ay6/GbM2dPlh0waRbpUvwLoqOB
NHhUQu5NoXwOnynMFutsCFPsyqkxauDKvV1a86oyendE0IFiOnjY3q13KoVEQ9czb9XW8eqzpiPh
zaV4WNccMZEsBTKjJ4JYcVvv6xTgzLQZQswjM8q3vnGOrXfFwOAv5M3sGKVcvSn2puyVxjYMptyT
MJLOTeUVBSW5JxU5soPoTBu5KYNGVNa6NQW8ivLUMDBOooFZJFqM0eZcoela1Ab0h4tRQeqSjlzZ
To3CYMBP9IF3a/KRK6xiJX75dV076fBy+4OSOytzaBp/kRxWDSWp1NZnxUniuP4y2zNusshJOkWp
lL/I+trVSJsTMuwSvt6NoQNl7DiJMTrnzHNgk5rfYSkX0emyrPx/BeHQ1oeb9cUCt0AK5vuUUauV
uWbr+ZAX61VH1gcVI0yhR/85/iVm0CWewbfXnBohO+4mRlcY6IYuqk7LBdsmBx6jFbGw//fq2qie
eaGXq6AQjDXJGZWVwUJPHIz2vVACpsV50bWPrdkXpOdXkGrRqOpASoWeW0Req++RhZ4nZ3n1c0vC
wZ6BT0AC+3IhturRfSBZbK1XSvWY0Lnq7w/+wogqYak+FLmon2gnV2ThJ3ju3aYP/WxQsQeByi9B
YwCEub8yCDeYSmlMvkMJ4Dzo+BGjbdNntUlZdUSrpTOrr/Studyqq0cncfPlx3NjjFoXvHwbPBxW
pC8muLpuyS0do4QHwzHrhVFJVkM3ruzBJIweqvA5FWQ8wJlOXEbaJk5VVzUh6/acTcNU1QZSaqi3
KifbNiDKJVFCxV9f70n4eJRrkYPjoNF/gi3E/lqsiIHMVe13I6wd1ZqqXnfPpaZyLnPtGWrHU/Ao
vD1bgf65NcZbTubMZR2ZP8GlHOJhzVzIIP+lUzdobok0scaWQSaFr78z4x0Ro/5Yqt1Ui6kzY5DC
CDrLZMlxt6S6XeGwvcB+fTrH7ipx5R3XFP6h2/PEq2Hb3Ex0Rx4hp5i4ah/tF4LGDkvKC79qblGE
qFczFd/edqmfIwHx6N3w1MjtRJO0KUSfhF9eRyTp44qWq45hjZVZN46OuypXTrVAdrmtka6FhG29
jTk+SArMsvcdW4u6wcNHrHNvq4FhLgicy+I5vW8ObAeQ9RxF7im/u8j2TNUPfHOU+FD9wBXALbKP
DIdWmcpUt6HP3owpyUnbLiof4+0ucft70YMq7cPqisMHMQTPlUBhb93ELXTr4/Ww27CbIWGhMqJR
xZbRMURdnZGJwE/E3JTDECyq0mwMUthvNED5tIW8hCZ0nxHVlWqcFHe+L0xGt9IO4hHSu9kRBigh
+jXAQijhi2JAO+7D46Bg3J6o17w4+UwAo3cSbSHqtuNDswLbCTC/lN5CJCk22ojcrDS/6Ep+hSxe
NSFKGTaB8hj10/Ksm7Yyv7jCrr2LoQz/NrRSyy7gwvnds+kng2TMRoUL7LbipUwA2WAzcFvtVwUE
4zu8UfIg/ka69XGAaJy79Fm/DOu82sixpmD9aFGJXFZMWuU685lZLMnuZ2UuzUj/PgwLbm+8m+eE
wrTve2YVj2jVVjXASIR3Z0Xt39Ra+G5SKYwddCkkCSVBYxZJ/SJR/cm4nOQJKYizsqATpc5rmlWG
f0N4ieXkZAE5IgczyZqfov2UH0qY5oDxn00K1eqjHvqHY4OqNJcKYAfbUSq9GctEen0P6ZULL9X9
cpytHRJbZaShanTMS7OxcE3PNLo0aqSqwdLshOj9UDoDp1SOJkEJumXejdsbnUPN6iZvqEAu3jNK
HgPpEvh1u9716OjtoChgH9DVMAEcEQHP9vbA82TVzNmop4hXD7I9oVti5WEIE1Gg1fpHtLtrsEUx
+iHRkhEYu6cnzO79jSTnfYxqCtEes4s9KH9rfxn8qiBoblka6/Y9HNNVMUuTfeyEJdj1g91IJWHK
WlDP/Xt950OOanbSl/KkP/s5ew2NZomRQvXgzDzVS6lJFDD0vUr4yRLFUZZCa7UNlgCUGdCMFcF0
LcHN6Crdghmnp7o+Yfnvb1Xen1zT15fHGVkFI1/ihRgkUCuH3IDDOZ8GsEzw9JFF2lFmX+YWnMZn
3Pr0ieT6UjLpcG27X1TFUwP4wwLnNB0Fw84vBIPtqwAEf7i+vQlYCWtNRTMmCXxki6IFwQNKkswf
/Q4eLTsqjePpFprl9Nf2fPQRWwjFeDjGgbn4WxkF+vFU/vs8cuu096e7IuqXNG8MRRiUH/8tzfSh
Q62Adclzo7yiLqAEyon7e2n4FXP0NLQMYlIajNjVtDUfMdj9lBibMC16M0rRp3EOT/y9tce2SS1c
Mg9VPJ/wcDcJlL862yOoYBFtbuVU1xSlgEjGfXPgekBqOPOW8kYQvFtYtIW9UEgJtxVEEWh5vKi/
mk2CObkhJJe3dcCusc0L/0oCVGep0GoInboz8TRkZm71WRSsZGxV9xGRdQo6RcJQIkprYiPKdqr/
2jsVXhUbAhu5vFD0tGtqqF6YQ2GAskovorBEQ1mFRxta4Tx4nqVX5X0Er7VQeSmRWXn3iM/M+wrQ
zZf/y8HCmcFWjpfChGQ/CDPgqAu9eeHr05FMpKKqj7Y+j7UbWNWnyl/4BABMAkJwRl4pwOqGYaqk
I/6mQNXVcD7xNaZiIDHenC6PeOKcohzQwa76FGuv+Pu5rMnWAskF9rNJvDpve8kXUBG0BY2sXPW/
YZ5of4AKHG5M3AvRdqn0pnDmYlNgo8wfk4GyX8skW3syVkXcPdEjyLKkZUgjxJJJcBnXH35PUR1s
11w0apu8zT+pmjnfkfEHreskxferHomoMRyutfczboS8GPfIm0zY6A5+OzWgL0+0hXbrAmxN2qSg
QNV9Ooi8G79/kGi3GCXRsxptUlWp9BN5SZKNawKbusPpxvFE9+5sD45tKQMwpb9gjci/cWJtHnIQ
F+eEmCHDGZavdMIqlX00sQ9EP23IjtMQaJabLcQke2i1ozW/+CBNw1FQ3qHloNjB8NaNTsf3lj2Z
TU8mfizxMqkH1CNvCShVbLtTKIRxgPAFZuDXKZXjz0X66TDFjhrQfb5k1BXEGuS75Bt64v91JkOo
+Cgme/H5pB5Xq2Ent8ay1mKZvFTya9h37jNCqT+dNy4Jx+Bgw1ag4n+5a4psCwKsB8DxBTHzs/an
1F5yFokk+rYtJlKgh5EXLeGtP3psOwwfAobl9YcME1jDzqAtJfJ2LSH4nA1MP//USTXNaP/5eSWa
XwXEiRFq2teDbBw0n2vNklkO1bf+l/YXW/lXNXkQQoqjAPyzOwvpSnpIz9hovhPUNClqiUo8eHDv
Fh5foLOqL3fa52SghGFY4Dp3Dx3a615FNbbrwdC+WPIonPu9n7s9ZPq9cRdowUQewEYO7PuV+cn/
TZx7ZzW3Brtc1j5U68HieYKLZEuJAr0ob848+3Q3DMFHL/x2GIniMRFeFnOaTBVXRQ+wlFqCE8us
9eEGKS+Y9Oz9VOtC94pRJQ4zgY2Hhk+21FWjcmcUR1csQhuLJc8ZGi6vknnA8qvdOu/0nnt0SciP
lGOxvRlaI5gPFUqhlBy5HlFh8nmjqpDGvjIL67ITAkxBxnUyB+dhePZG8JjThhzYyplo7IOxUlXZ
ROTKdEtGz2j6dnzfOSvD6d47/DNmBkaShaPMIjLC6KR0TWKRWZ/Jl8tQrnYBkK1xBX5gw4LFTMZJ
QG8kQxidGMvLwCajUhqr8ILBUktA1YMIWrNEQiJ16A6Vbfsph8KcPfb2LM7Vp5YvhCzIRJ31iH4W
P69hGCO2V4mGLzvNW8S7LHGwbeCx0ntwijGa1AF7h/fJB3hywobFiFI1gGwzSk7h1ya0b8ZgwsMW
a/xPpnyQXmkKvWUSpUzKOSGDhr3V0TnkLeOFRACPwe8Sx96kB6889pPwjyWIlypqtcTPOrMfc/jB
uHd6jKjCFd9bG+Z6c/CC4j53UP1Uw2WLuOpni5zcKxdNxwXNZATf+bgQOjC8ikhhM2Zf5z3Gi6KY
0I/dcaM1uMNF+Cw0zQ7Y7MrxIIR7j8eCMJ2ijPRwnfsGi0WzVk1bWoGMsLK5/R2Lsi9igLgLN7uI
wT1mqx8JmIklcHz/BTowNV4+hJFPAeyhMRNcZUdEhaTM8pkdXQ8fZS3Olry6nwg7jC6PLCxwz8P8
KbmLm/94F8s0QY6iw/I5Vj0z2hRvTDpiNvxGJbH1FHlhHs16L7a5WHw7VCyKu7LYl8RfXP06yl+c
vG6moJ/MZsIkEXl89fknK50OGMAa8o3p7oJggkEaxkHxgnsU0kswgvbfaX3e8+7eobBryy/DFhex
hrxFLgp8Xm8/R6UjtRAPHe5UTmbkMfnDG0+lk9J4li+pa8WwnQgIidxlX1uJ+lSeyQwyWjTw/8Jj
C77+vTRdk/txMVF2fjEDwW4LPOadpUYDE8X1KpDz5cZ2BR1DhbWFkwtlrYa/F9JaohdphWONt2fj
zUHMOoRBHiTux12d1MG24CoDFq078Ip8gn9FdAqr7EnoqckO7Pm07UKESl/Zplg9MuXvdddsjRqU
JQ5U9LoBt+qOS38FJLkrV7pwYfugmsTdoTrPBPpYE16IDsWxkCoUSKY+xfYZROr+AsVT1s6T7Ky2
Zf2OQs4LUVB09zw+oggD1OWPp/0ZU1f/QzaOK9Bts+lGyhO84jKPwmR+Q+jbhLXRJuCWjYq2Brs6
V3vobz9diXaVYEzdPaEgAh6oKx1Z+1DNgndJ2PZAYvofXSyttgFiJbEgl6mr7WQcTUDp5/1aDMOC
qZYs2s2dFGvB1DM3fXthlwxr04zCGxjvT/ksNAK85aW5btjus2StGR7o27euOJUKdwy3DrjbnlzH
xacyqhMMiH2tT8CTY2uhOtzWJ8+P7WvKVmwBGy+8K/er9GAEXaZ6t1yF66oO7qNjkUxcymbkZY1T
AXay7KL7I/Nm8U4LVzlUMNZEnWCkTV8tkscK8i1W7MiP5qrsiYa5jZT+XpG6VxJyzrnozc1Yoeaz
QH8Smv8n8Km5snlLV9otEHSCWPgcoIzHIW8pliduiEwy/P7UURKGxSvLxWRb61D7RwVoLblYIJd1
e80+xRqV+/g2gV8eH4ZX1KdeemoaWIzyNY3i5KVgS0tPGrxvDkv1N5o9aREgUg6nTqmWGsuDocM2
T/6UkFlv822kvhvy96gNK9Kk/OJ+OStnnI4o5WZA6DjTc2Vw631vtQD5MjCRuF7wRYK39LXevXY0
TISM6dQ3QrtB/xjhZZ+FJbfvrXHtJphuGuctRqsvPi32e93eddFbRQONzSKp9NCqhH242rqYzCk9
RlFsEJpvAlxYCeECIm0bh19Dp03LAk+2qWN+XvxpkYTnmRv9M2UBJalpNlBo3PNcaf/kbbMhHnuk
N8i2jyAfCBVQGc8FiIoCH30vfTMnrnoonrHXfPG7Dx6jba87hH+DEq9sKpQ0bwNKF2Rmn5IKcJVj
GmfzKx8o0LfKCedOA5ygbgWyWGcJJ7yeR73ZWDRQMd/7CXw/Vsfq6sH2YHHQZ9c92ciEtIApIEUr
lEcUwG6v8z3fxbcxeiifbL04/MpK4Kaqcfx0uI2qK0wflswJge1jn3mS8ZLao+gzV5h1pXv8YxJj
Zoh/fLGUWGlp/UlGd328O49EZd2VLyJ2bA6iLa9zqbh4ZKOFi0AuokjTCYSbZQAiDMOsTnt9CFBZ
VA5Kw75CaCSzcv1V7rc6LNxFfQ5OvIuUS3DUPJkILNJV8TRxNyMddXNARDoHqQw7uHtufM+kZwxN
Wz3uMhfJInsGo1mwOiD55TKs7mVvwNh3ocTAVOr1dcBvNwOhtpeKDSqF/QHVm0jcv6rfmW4zusS4
qWTElTcBrjV0ZqRcgokDyZH2u4dHQhOmi7KQ4dogBLeeK4kYTWteMjTA/2pE8CSpyIhFJwbIxoRj
H7YzYCkO68MY7mBRJJbeF+YWTJP5+gpm20pSV7xP0fwpKHbcFuVVTX6YRtEcTrV258V5YQzPNaCQ
Nw78JGyJyvUiCzRk2AwWEA4ndYzKZhuIlgnvzc9Mx3i/Dna8CKV7V3wpd564oi/RxAOVvebvXsnp
2fR6VRqD8iq4YVyvAon1lQdWpBFuDrUHcwx7K8+H2Auc0giCPI/ZWhr42k3aKI1jv3sowIxmeRgQ
iDxP4KCM5lb+V0eNZw3KLVmtCJ75gboRA6Fx8aA/gN/Q9cUJK71brsC96ddZCRBQv/fh6Pv34+EA
+Wh+3aHRtdITRdg9ZQDMf1vbk5tcagLOi8YNhc2gFFgs4cz8tumRut79z1F8Fh8xmOVGxOliypWi
JWCKlrG0O5cmHEttkLDa6Y4+3v7jHKljM07alx+4ACZfCnP4duava+ZhVYAwUQvSjZ5pxwfacNsT
G1mMSXhCNL3neIYXFnWuvbxw6gyVo7Tk98LAqW8XwIv6PUfh6TBSsNZ1REWZjaQYXJFpd6mHTHI2
ih+VPOtFIAaGqDAYUFaGs4s9hszxOwTc1jjQl3kQ+58g8mqH79cGm+lpKmJGxSMyh8epooVwws5J
EhCC45zq9F73FbDzUqHYKK7m3ChSLHFW+dgHQ3sYTKs+iF21KAAD6iEZtJ8t8FHTFKZCWD/btR2X
2enVQtGFK6dl8cURthbR0s0xcdPcZUtE6P27E/1WNhl1DnQf9tDFvrP3mVKNaClZFBvF/oFQp9Fo
xU8i0revDP4mFwlF9s3GDnb8mJQSAbO9/+VwNGsfdJkKtits3m7adqXwIRMJ47JTY2ufxJGCyvSb
yNm+jNMg0nxRtufnbvfEu0BSUwzWpzekMczbBiYSxPYnW+5NHrdCPP6fvMELBaxuv4USH1EkHbAf
5aMu3w+S7AEN1kF0920lBunp9MgaVdvzzV+hYePDJ/mSxH5rkvMoBJQAY69ebV5eVLxVnnsQsTaz
Qy8DWN8gIZbDOCkGSZMGkpn7MO7gGYf4atJulc6wNOH31DbsUH6UyynY1J9YOWErkz+eIZzV+Ep4
igKvZ/esvhM0MIELn7m7Ojs+8cl1xH7JGnHizcnb9nBG1Zum4Wg+NB9Cr7S8AYptsfI1xImDRg3c
StgTJccsa8+vTF0FIKLs20mq8SXYP7fgcRe7CAViwxfsLokkw0dLaAoKPk76vz/RLRiGICrxlf9r
52AO+NxEKuNLLMkmmil+OdHpWLcEz6bRsHZPuVEuuuaDV936oA0CIGgqDUStuBlrsIzxuq10DJ+F
iTx+E0j6FzaEa9XgJH2eKUomrhd0mgu9QbDhYjjKFGC4OXSlGpd+KNk1bcUsTcIv9XgIs2OGYQ3I
Oz6zhlBwEk5KSNpt2BN9quM6Z7g1zohGYVmRA3C+DFXC+F+pxsauJib4SnHfDHkrMuQHLlJ4qH/k
iEfHabjC52TsJFT1cvWNh0AjRlRyGzToVvT+67OeMrKT7ud7wCdqOhZBEi/2e2AxTecqGjcdyont
kE0QamkCw2ZWK3Eu2X0jiT9uezs3Jq+NQN2t5T3rncz3e4Fb7KGhCAiENFeXHHpQl1DN6W8SWbeg
2AIuTC8YTbanX9BR+Z5ZEsIbLLL9YCs/N3NFimejIz9UvgVI0HLTl7p62U5xqJdkFn0u7cyrQ6TC
bElFGehsZDKAFOWf8ZsldIBO3TcEyTf2QkuWismSSpGKtmJYYaS7oEZ7V0ydSWBA4LZoOLQTKqbx
8b5tXmd3N9yt18GYVrMb6Nr7BNzW8p9yDIO3QQhOPcL92HM0rQpridI268Q8wXkp/E6EUJFy02Lv
tMWie9qWKAJcyWdZNuUeTi2KjQUk7/6WPSKnMeDJk5eWMtQv7Pou8zH0Fv/5EuD7wt3S5ICm9l21
w9bf5h0vnUsOg2tlNIh5h2iu3hH82f6qP5Z5hWUR+or+UhDxvlCMl5nqqdvK+gounXxZR82O5rxH
XdowUSE5/IF+aaDe+EIDphrD3azfOxUDFArRPN77fXSinWRxrapmt3HXZpnvXlr5oFv14MMaNX+4
Uo3zso/c2JlUcPKlxF3uSuhmWh1IUPqppBnhjL07Y75y62EJTaz15S0F+9MTB/ha3keeR6RnXUOc
uwIENE5CSRPurRygxq+PXWvhT7+pvPs50i+m1ETxi9rd/55COOQkaIPdbN2Wm6Je2R3ZPH7ANPWR
4KsiZo4J4xriEAh+v/9rkaIbcATO4L/dd/tDCIP1uanMGEN/LDkIC/4LSwZwCC28Ni+foDzz2vnv
/vslzLXLCaATJaQ+rxiMsYIJAguIgSikfY+adOvLU4xM4Ao+pIj+6Vj1jPKLPyqlKIcWhcMwskYc
s6QR3f8pw95nGi0UkOMle35WCunqFhI4EKbGkkEfj3GALJFu5YzHPXyz9oJ1s4iCkMc4Hf1yN+KZ
V9m1BoI4LD4MAFszW1bmI7uungV+xLG392k7X0LY2L7TSO0AP16Zj1gKv4cPk0qvHq9TIMcjNxJQ
83mvFk3L1j99idDb+rw7dvjN6h00S+mXpTzCQauERFV2nelHFYSLENPOf8wCLrU4eSZKyjFrg9I7
uX/bUaiZV6B6lamFMdOJU7pTva2l4Zwvh0d3RYJuImWypLFtVhfB+yG2VG6sCTmFPczkwaqbb/1D
TY8kIFfXpGKvwrJ41XUt8haVd+FpqYCCOM7hcMI/n+P4rxrBh3Pqc/RVZoDy2ggglSRLdCG0iki8
w3Kmy9grTNq56ttYl0A3OwMwA1LV8f2ytMHzSE38NaVQqIXzEyT3HNFxhz8NdsWtj6s9+1w5Op7u
MDa5+f+x2x0D6esG6KAXCnYGDYQ+JvzF2xDdi3MnqCJ6HgnD27Q6l7TqHj0zmYZvTFZ5oFghfdcH
pDmgoIbYs606UiUW+7VKTENCj7eiH1dfXu6jsqv8bealOmabzVtpxC8e9wiEZkeu2zIvilIeiV0x
B3a8J4OjLL/ZnrPr5K4AQ1/bBWTvldq4XjZvYTYxFk4zEp46hzK8qzdDkgqtESwZp63ZbojDvrdo
ViPFSNpRMgLUtFfBQZQB9DXKbmD68V9GWemHPT+UFZZd9PDXhFQiCkg6im8JDlYj0nQWaQ68k97U
LO0x6cPgTzgm+qUsdBw8GkTtTm/1q7am3kXL2jqRcaQwYpSQhTtprrzOaCyUhUYJ/CVanw9l2dMj
PGSWlswaQftM73vDFVASVTJEkZ8Ttj6d0IGiE+uKVdBuMlDCvs03ONpkgroFs4XEedEMJpnggbe3
a6PiW9V3HWJvtKCYstQ3lqEWotjZhaJWWorQJLG9ztuuPnu9wNsIUoIwX5bAKsF5O7tLfSEs5G+m
y+09LhBzfx4fYyNFLeNhGB1ksAqLOX/clXJzsEUs5aY2yuTUzQCy1cLY6GC4sOAIjrjYAX/bW12K
VOycuyL4zCUyXlI2x7m4sX1Zg4UTge9GUEIRLFmyeC0x2TQZjWoiZP4Ez6QYwq0h5dM21JfcGidG
0+D/mVBgcvHWAJTiT8QxyRDhaCfyS4k+FfAxS4/OZQN2PyEt94ZLYtEZ4itjwMmY5FqQWwi13hW3
teWrVy4IwXF1YVikxnpIOJdxN8q8cauIp6Jh7+Meet2LCxufkO/xUaN9kfE99+nw+7lnc3s5QyYb
f0yLPceBUCGQkbouxIjoB+yGZE9qA/Mg3HD5BgSD4e3ScFm7bJ/lF+XoF2R1cLIxi60nHV5Y/3H+
SxNZpyz2o60JXIc/JFWn9rSK9E+8cQaWKn/yKyT3BZSwKsKwjUWixtw7NiySho0KCWL4BmB3QapW
3cDtnyz06NyXJ63P9R2120jFFTcX1KyqI5gm3Xc+clf/Yy3BOYo2ORARg03YarLPh6u69fgwrZRj
BKT6lGw8gGnLzAMZ5B4b4gBe1Loh1DR9rYQhtMl2y6HJscGcsNWD57rpIphw0u/VSK5hRGcmaxZF
/2aTohktF6Sr3SsgeATNgKVMqcLTmqyodcR2F70bRn7r67K2wUO+hcxwxJaLA0KDIrTkOPmkCxMd
7CGNKou+9HgQFzfw26YsUeIqywachSZB+iwq/6ASfWhgirXP8+CpzrWGhhGIbckk0BYuo8s2TzZE
DCJCTumBHHmdki89PHxgmHt1iXTCYkpfus+XWNhReujBNZ1DbJd/BB39MoIJLRMskVIMkQsnpxHd
RFLS8Uvs4TRcXBfSrzmVm4b83MrMEj7R5aDU/NMsfUCbn2I564h2ZAeqwnupXww+ddKh53TINKDk
PmFpurzBo97MYZTURs3m8nZWtgooyCTz2raKI5rybHz3SwJFfl+YM2mLMRtXDOL+qVojVcQT+ePo
HTbhrCYOq5t8Sjuy/BLoec8E2i9ihQMrl/KehQYK7jP+7aUenUaKw3Up8xrChS876Kuj/K7U5ggB
FHtMQdkc+4W2u9J2hMyRtpcN391pvsAedTHvojMOmAwPDvepwJGIVCtqWSv9OMxfW44X/0MbKsYY
OjhCR+4g1TZU5PyXeGEejyMWJaIxGv/5dXLyYvRJ/znSW4/c2OB2uqVJZUSx0DWf55EOydQ7jwwK
t/fDmkI1s0vB+h4fZzG7/GVy1otc6a8Cxi71PNTdmkqr0RJJ+vs1cR9U0Sy5c+ZIwjfJ5/bvBRux
+aTdHenX6jyBkxg0ZiVi+21ID5bb824MCRmB/gfLAz1gHgePLvDOJi/vQzVwRIQNZJ11wVR9t5gg
I1PSgklJSid19eypoFY328TSdcIhN8WDIFWfoA+YsjSXYql4z7EAuLj8W3u9oinTre9jTEWG0uyH
QA6X8OxMuXxPsuLNPWYSgTYyO8+6AncMTYLpjk6VoOHyuk5JsHRGBtxRxFIwxJYg5DAQGWIXi5YX
L0kHUM0Ye2APB53Io9FRE4aIOSbzsGQWZRnFAqBBgqXJ/lCsCTdxqJcYOGJmOORP529mVyUo3x5W
P4wt8T7The/BHTnx8YNPBaLJVCJQezzrhnJ633f645QwbwJmqAv5LPk4GYOOFxJLxyM/+hEOFtHU
gTf6IK01oWEwIqEXa3Yj/t7UjnLViDEasecg6F5xWeDzWrGwgu2icfxIPWXR0OLCEPAfhvSb4YTY
6ndM2teugI3avwGi8PD/erNn30jst1Hg5IyYBTJ6YJeWBOVr/wLJOM9DOmmgLEQ1+NBU06ZfwpWv
LmUbA/jo5SUltr8h58vj1cgUHR9w/jP3ZCiu87kewc6YnaUFAleulqDXDabpLX1NiWOrCybm1IxJ
69BkpASn0j47+tE6OxxnykjDU/Ll93DN5SbQGxbD2+dlkaelFYT3DJ2zo6ZTN5B0v1SAyM5OVY90
tbbZnrlVRig0/mtD9l+ksW5dXEj5WaJd7fKMQfhVBqhovJ5lSZRWaswhsDO1Tgt/YDCcNvTXgNmt
+0jAg/HxIX28tygoXNBiQ0hZ3QrsgY7hvk0bp7+dfuRn3cWCnWDwF3zNitChmhsQDLCJrCFAmVjf
Pe+cJaRRf/S2vyuXYoUhT47q6GQ83hYs/xz2C3158oLYgC6rTDHKIjOpVUAq1q4Km57Ms6f0R2jp
kNInL85qChKdHdFBfTf5pJiTEfSfG7Tdmsnb16cJRCbOJoEazjxKitLf9Xzp9SWkR8pkObfnoVBa
25sjMVZBApbjAmCVdkkKSoIRc3A7Td6eAgjx7PE/OExWYk0Wojup5xnAgLYsoElc2kcgA1mpr4Dd
FrNxpHcXCZ42cchOJOsex4PQkW1PdqbLqfsXvZMxXthpTl2+Vr8Kxnk3KY88zR+WfTCtLGTK2NqW
IxvmKp9SlSrjZCpMgdnQ3Zol8BOhZWAZb/YIpZgCeVEGcTviKXjE451vW8ygMLXDd0Tiw3wKZ6m1
aD9Utc2ZzUZkgvZvsJzmqpJx2C0q6d5RFDVj0Uwxku+9uy563XmrXdi9IT4pw8EembX+kuOVrfNx
8WxBZtj5PnI8zcYmWWbagMBX/mgWe7e0q68iIaq6ioD8XfflYJCLwQcnluAYudBs8uJn4PcFSuKg
He3FptEWY1B+CakK4z9NWnPLcmLUHfHpzuPS36PHAExPBW80r/u3T+4z3H394XN1bV1+ZCcje8fA
9JOpeb53hk0Nq3xsjUmJ+kr+Q9llgYqwCjFDM4tdMOkpPgs+NNDUGBvnP+SfcD7FcfFmHGiTMMSw
+e2OdctlYoaxh7sekew6bGpa0n4e56UNH/qkBQ5FOmi7mPjHzmfjzS0JCEd3JMxjPihvXXXqTbjb
hM04xjtgbo0yKFJqsRiMrjHA44sHTOk9U5CSU7TjDL3NYT8JDz/1FDCNBr7DX6w8LPuOHdOmG9p6
yD92oH2l4lbzdK8n+ayo06sA35MhJAQstnh36Im0gfg2EazZ4ZcR+brabTH2G/A8bbSiK8JB3WSX
P67Z4mwSzEAImqawgBCcQzbWsnoNxsTw8Nedv1+8edOl+S0ZPdTcNI6cadOnG1P7sFJTnecIPouL
hZl2Fi1iQJhyxXOilLMjiiXr12emECWj5yBgGZnYPXpR0nP7jdKNfYpsxnuQG0ywxn+/r0yEsu6T
6xWPvPPG0p/y4wY0KmCvpGS8EK70HBsnSHs9uTXJRncACFfIR7lasipUrmB0NPUCtaOWuzWNBHFH
VCYqTwZNANj36KUSHM8rY5yscyOpoBXZ0wEinkBdb+t90Oi7HXQ83uDdU0LrrdvuBg04u+k/9Ehz
qIsC72Dms8u4j7QIGmnohAJdtGqQyqRuxlDFRmxK8FChUfyu5zWtPF3AjKceBuf8UaUuU5BUkn39
n5Cb4xmq2NtDjrMvSTgUmMadEQkdYZxZeLKUskLvCuN6YyZdt85l2dNQg3moHl8/e6dLIS2xhVAJ
B+qdKLIxjRyzzAgphMYM0yCyJOgmK0ca2e32kf/7EhYdZlJloLqYdz8sk/fSi6mAwg4ct1wSECIf
9APBGWtqPQPLn8DC/FLvURkOTaRQonQo4wT44gtUFsFCBqJiBnTjxm0ppGjMyNC7N7k1EwkRZg9p
5tfpjdkd6KfrMw4iwMgEu+NMciSOpxnSKLOiVBrBPMnGhduzCps91Bs4eK5rYrJ7Qcewfglgdrre
EpDV6otQSeKWtEYvtZq44dFP5spky1gQ2MzDBfYq7nqcNfVehXmpSA5nmsxOCQGEzEH6EVZSAMl4
gpCcmof3c8QvE40f5YeogXMgso9UUmInbntqvBCn3x0uikQ2MSSxHCT/oOvxPO2/kwmW5utk5CxH
RbXIXLd4mYji9xI5m1yEnQhPSsq4p5cXFWKYuc/bZAREdGhfZpUc/qA5mIID9St84AlBDbzOUhqT
Bi17/obAp+u3F8WgiN/KD7nfaIbU5TctqppfmVxRozc81KNRvN3caHeUzlxeGqEblfQ6ban1lXnc
LPHnh+Q2BurGD8d1WG2jABSEcvaVKSalDOaqUAySpvQA8oLoIribpeMmOe/OaZuHGdnSCCdzwIdd
Gpmg4hgFDbwIJWs5LEh70kPGPc4VKNEOQYRh3ug2x95feXIhAqD51Jbg9aF+y9bg96QQlDdPF3Jm
rLWXKyr5g9+uuKuLBZXnss42YWSliTQupgBiMuFLKxE8NikYe8HEcCQH76rSIEq4fUzldDhUR4Np
EpLUOlVqkLLD42vDf+leK6rNgyCpQ+/yWlV1nmpbWPSU4qNpG0HNDVvaSy4ovqvPCs31NiZQxScl
lDF4qYQyM6BtPsYzwp50FBeMHMYffUZbk9C8uev2N8wLwMz/Mi+fv7BKPE/lq882+F80dCP3QpxY
Vu76HbTpL6QVKGqIflhgL+OJjrp1OGgeXFt9P0nfgo8+z9DF54uVdi+ZVlEwkO2vXS94LVRsUnfR
rOlBFm0qzzhTUfzBOVdi8539C7JAfwUoSr9C3bUScqQ8VHrhsGr6VITqOMyVeqE9CEJfH8MAlnmu
M3JXM6KfAw+QS65GZJsJHWStQYrAwF+HF//hXnJTDEqYHu7OvyPLnIZf6hyU1ows/0Px+2ezlwWU
te9uHto7X8XpxCAd5CT2c5CHiO7JS5+VQ+0bOavNH5w2/0Xh2+LdD6E3VXd9MorpCmwrVPlZmvRn
xAELTN/WdFQgQOvHzUy/IGcVVQaqP//aSR4saff3b6SfUwWlA5IBooYaUTB2yLr3pxONoZrIkVTY
K0S/g60LENzKUvXFEe/MbVx2zBFkxTyAKgS29fjN77RWp4tEO13KwyHRVdLpw+iiWbkBZmczTgR+
BZRMIOBqpSuW1D2HBDNCbWBW9G2q83ukFd2NXTdWZ7eJf2NMvM/4mk2LMJcRn5tKJLFuA2st0ROU
1kqH1OgVvN4I/eEGO7YVI6QsyQ7QYrgzfTEZL8kh/Ok21QypJVzmOVOEvHV0H+QdI3gO8bIz7ovD
xQc3Y2Y9g8R/RqMWBffhv+iqi+IeG7/Ai1TKcHh2nvZ/ZoAQAW/68oj6OgGteQZ81ZAMCGPU4vIl
cqYAfJGkI78EaaN5oUlll9KrPbCiRzTOzTnMYyOFxyv7O73DDxJ0/VjZKOFkDUgOJfpA+jLwX3uy
B2DHDbvIUOAgVOW7vsIjDYuttKzQWctw1l2Rl/t4K3ELdf5SjLwqqaz0nbj/WT/rjiZb+KZmRq7d
rtUqDr/HFq3KgrCVMGOz0PgTelGc3FQvMe6UvqfoFR77ACHYAt8zvT5UAdYs9UcxLasqfmqkzdAJ
x1spPtar8iy3Dh7TYAd3qEgcHkJUxDK3hEU9nSCn49lAu/rX8t862dyn3u7tsFVfRWQ+G3zUp55E
8NOf3GZ4nLCvCbTdE+S6OKzJKKdLXCHCmBdyL/wqOw5KpfNAWQQPkeB6uAbe5s5piWwC6huk+4EL
tCvnnqii6iDhVYkp5/w1xHaOCVsHtYRie/Z4mO2WJaP5wdN63kSDOMbexRhk8msgKjnD89TDuIys
zTj92+BrbMuVN6Q5anfU4KcwC9tGkdkAF6vi2oIqqHactL/kSpt7x96/X92bLpiitUsJcoSB/xWj
HwEhIEtBwO+VwcNr4FNW8IX88Xf/op9HQLqOtvRv4V2tSPIEscpW1j8T1KNLrF0dVUWTTsWAJL4T
4olviAWkmIq6CEABtn+7oOvao6Z+nA8Oe9v3KhwbduWBZHrSy/ZwloqMqO8uN38wyyvEAi1xh4fz
BwwQvh3Dqawky1XUX9SfCSWOvEi8jAmFwX5hR9zNIcEI06iD0rXLCgVnfXzX3g/zZk7EGcHEq4bg
blNLwLRdPKJYpoujUnTaOP5EHFldP5+h/54bUfLVKMfwUfSiRAaTorIaB6n3ZvRyhFG4rCkdrdTJ
O72Y/CP8ocYoQTwvYM3x7t9oVJ4nrvqFvb7oZfYIEcrcj8mZ4iLiLmviqAceQBFpfa/OjK/rPpfv
5/SSj/81WJJf1SKsFoTjA7LAebohXOqpKc3QliXPdUeY+JuXMelZGPgpwWcM9PHQNBi6f0OAQr7d
OCZ5Wosw93CUyEJ2tjqu2Ap2mgKq9QKxNf4VREzoc1Yr396AI7cJHu8TvIBCzT0umeonrrHVJ8fZ
JweJum6orxoTQt7TB+2PcO77qSTAGVecb1MmcPR7TU07y/cLlHi0JFKevClpFNEIKBL2RBq7LMA9
BIdvCHFVzLXF7DzVSZTqXNkJkG1vo/clyupap076cVcK5ZPqPB+eL0OrLoLONYVHbX8UNXobz01d
DHq8BwgCbkXRZNwlbCinrpM+BKPgDFLozip+yI95uB10sPhFTIWi+n2p52vW1ParQXr/XzWIdb55
VDiwxJc+RppBVjK2QpLFZSRIA5AszTIipbQU8SQDm0vdLm5Q5ehv7AF/REph+ZVp9IhExRKzh2V/
Yc5oDSSGmCGDp9WSZV+ueaiEh4KlGoq3gf6IA6dUjie7HwZfH2j8/YBF+Bd9IFMNwDJN/9UA4Ciz
UBvNfIW+fCLntwEaghLIJkEtSUZyBNrUKUGtVsrn0i3q+K1qfFf+tWjGjGh7kfsz/xgpjEBE0fhL
Y5YFczGYe6VklERTJ7QdGD6BcBaAn2HNH0uNFuMuMW1OQ9tO/n2eGl+zutC0/Iv2Doe1481zCQsI
1jSaEpD66KSi25sOFcEgevOcfGS3Fy/TwtYoK0JexBiViIcW9xIKWGUjuah4+k3/7yHq68Axw8Dc
PPs6R89axJjrwpmhC3WPtwaLYKw39RD4emz5Hl7ErIEf8mwaW824AH+9DzpTKD2iVUWr7ZBV4Euc
6vsgOdYlLgWi7UKE17KFvUYQ9h9WY7qtXZP2OethxCC277PhLyt4x3VDkfrq/srMEsC+a/qN5kkO
ScYcS+qVCqVnd9OLWJ+f1wsA2iIU6NzADBluU5sz87w+TdkOuVF+dCPRLyoC8nXI+2CBLO+bOSVz
F2bdbgEx9YqF1wr1uflzHTQRyEiyDXRqp5wMDGlIGXhUEky2wiTV9j+D6VGvVICfZHzh0kb+IlGg
6XG9IkIrK9+JTfF+gEK2tcjSgnfYCsV4JDZew0IbOpWd9iHrS8G8cgf4jOlu5L9VRjnpry1t0Vil
kZCTBviPMYYmQxIUk5RvbhyK3cuimbWQY2TTvnwW0Se1DoDYIlyoeSzzvqqPxEMKX+1KJPp/nGjE
trGOHYqtp+S6HKIWLvRJ6lJXwbsw2qhayi9FuD8TeVe2QIuzAfAtllprX5VP1lyc8fxZsggFM//m
GK8PGk+n8f99jH+3vxTNpUVzIavPs7dWFUhjN89NaIpXRoZYnGj4bUJ9x5N+nyKdX9oiZf6Bx6Zu
ZzvD9jYB12Ab3qDgMwEnJQtMy7hA9MBj+K1cuFreCOYNnFBY7vj83NdfZca4F1eqNDMfZ2NLfpGS
t15DfY9seFvovp6c6QrEwD34kMw5TGKO0GqSZbtrRBBqyjHOBK5p8+lq5kU2lu2R5kT9ywrLJKDe
iueCLkD0dJDTKjIv62J26n96X5Xv6HS6ZQnTHYG7zjpnGfSjSFScmHWuoXwOFsXD+Rp2EsBYaXG+
TAg/rvolOYysNPK8uvZexyft64w/ueejUqNbrVIFaYZ8ghqTidVmjpE3/2l+R48emLeKpxtGzzuq
/1r1nYI9dZbJLGsEwzNtfYK7ibOzpUf6Fxp0C7NC8D0CAcR3YQNe/MqVtt//TDaQbwVsYlZBfHBD
G0NV0bZlJjZZFVmcI9vWEnoyMQCnHrIJs1EAFkdMTXNlsOaO8lPw3PsTnk+XWRaHPsL0HTTEnsiZ
Ye3CjKFrsIShz095snZZVouZb+OcjuFUJW6NKPHx4UyillqALhMZI7rK/f4LEVTBS5aEgCWUQjj/
n5aF/UL1I9wXB8cYCpVj6QGHDIQTUrJDrCfMGtpb7oMYL4LDDM0b4NUXSuAZDqU5g1Jujt+1HUPU
JbWhNnXFn4O+Y+Xx8n5W/K1TD+NpPEbisUlFk7xY8qCMqA3Ec0H893mb4r60bCc3ADwE4tUZjEsf
XQ7vxKoag+RRZPhG7GR0EFANcBoQwYuKuUYemHiI0nkQRvojYjb1vSDt9eNlb807GQKFwaGkJFcz
ZUCwyt06ThDTJPYOc5rrs3QBwck8jvxxMmB3+dAYkw9muACVXF6UBUmPmBE6CWW4771Y30aNFDrd
N0boxDh9EnafXKGJCOjQpTeB2jreAAP5ZTDgn5G5TiCmOcSkopRAraBktDkaZhsU5f1v2ba85am+
nks1bIye2jfxRmXaAdSmuZJGUJUU6OZinl1VHVtISNp+cCBo0nBWiHJrK5R2D8OIxkufYFJUJ4jm
miTmWEBAm/PV1YlMad85NbTnoAaNMRAh8tmHG3MCfVR/uT+lk2niEFuQUIiI+cfLpQMDWRrcwmt/
kUZ5x31K54BfRcMilS6A0swP5kWiXfjzPgBcy2Zw+NvEskYd4BIxKHzh0SKgUu+DCfQ37hiQoXfN
Ene7pbJvfWJbRLbN30yfmndv6fjy2XkNs45iEb0wmj/LAwDDeh8ZAOPdXks9cXYbGeFpc0YpKJtM
z8pUaH+051pbSUjobwmOBEOs48yvBC06/jvmL9iwo9HB9RwQyhHhnBpE2WVTV5ugH3N2Jj0nydBw
QPTN63XH5bOmOGa2CapCamgtwIK+YNyxfVzArFdvk0jC9T2fAwR3Jb/3ervvm8wZvBrbQwSUTLuy
NR3VAtEpYfiwH8Uc9fbbutbL9Ex+Q04a3V8LNxOImGFgSCEVGElcCdVicChrZwkLX4Z/FgrnSgaJ
Vm1KaPsEd655Gu7g/YQrMGOOL9zhqZQvQF0Dl2G0iIONpJ56WAVSnJeH/+xzmg7HsBcnwadCQcqW
wOlqUphOOqmpTGpA6FotF07/bgfXZepgaEPq6F8ADoQUZY/XpX9rari75nqNlxqDTJUyK8gr0tZA
Mh6RdpwcaJdPwvh42iALoApxH1VuNS867eUH9jmJjmPD/AXx3Rmq69SlIY9ghwpo1CfxNh4MDyIy
iBJtfEtMPPlJGXni/Jg/Y2rRbqFBuQuA1JBcgykMLfSGtStG0s2I8/1EnkLTESf8jfBbLxmlGMU+
C7rpUbPS2dCxa6wSqDwPIPlKKePGz8TfWP6xB77orpLS3wFBuC0wB1TJSKYqNwY0nK4s9yk5JI0X
FyGysRAJR/HTJfiAp8PJpz2+pDW2xlcKeeKmDHRYERQocrNBIBpR7lStDM3aTpElKX/sWEpwJbUr
yklC9+QLqZ11XwxSUgyNPKW2FfHfsbRstK3NrANd7kOplAuuU5okbQC7wEq2FHYiSNjLeyNPDu0W
lHzCaoL82oJweP+YcovCMiTUjwFb1V8gPu/9TQR2EVmv6O8EuyqwdnJfL7gpAmSE1Jiira83j5uo
J9PuDOVl/ejZJRjvwv0X1DTpY1g2hfrLMW+6mjFcPaUd0FBZcnRCiU6+o57h56uYE9zYEoWsPVjq
nMfH2/ZcxSpIP/salerCuQeKYV/zMZ5yReMFgFf1sLu4EWGvRUaALCA5KQ5RbByJYMOxL/qIKcZS
LNuLgoGszQG0xD9SW3IBq/1xBVw7+HKqU7/h++CINiun3n/ypJAkckxsp6MxcMH/cW0COeWyKNql
Kq1b+ZAF6YHt/IpbJDEt8WlRjJwsxQOfQnzbsbOuEvDCOYVhjPyytR38S3WV0Ct8m8W2AA+b9Akn
cjsBZrVsrmxEM7B8IPxNlrxvqF3B78fFqD0jVUhLUSj1WgZsxQjKX7PhYBPhJg64kmkzUeNAxRdV
AgnHbu5VSTZljfMyonl5zBmSOexTuPrHadZAn29sk2uB9wYTlKVNNu644ig4Ws4rgV/GiicHf2rI
0migySgykrHttfhDW7hwafAI3CKN/FsrDc4LmIeOjt8y8zd1XihsjdDckGDLqy/NQTGelSQZGT7i
vnXfcfPeU3VQAjGHj5NVadRu0sPpYWEmRyvUAyYN4VRE16n+w9a+poqE1rZ8/Mdill9CeXTSGO2q
n650roxDuoJpFTHxzOgdbHV063DRUarfQsDfz7Y8uYWmMLU8Ya8aorWusPLRC7LqJx8EOEQKWk07
h16fPWAH1WHvYqhhGawUkVzbF6YSp5ZXKo2ueTsocWNFPTZmD7V5kcNNRxhDMYDMLkULxxfFelng
FaKrKSX3XoQmT77dDh9deo/3dIEk5SG4nIjpLOIYOqA+UluI82pWiTWhLt6q9c0hbmV7PyiV8rZV
1uGelg7VU4kBVceRw+X4cHntSQOQiLm8NDZijCD4pXSC/dFhS/1W3kmYr7vxbv3oNQHLUz23LIBq
q6ZWWmw7x//6VJQLdpXNbMqFEokd6q0YTZgZrhpP7zFy9u7hHxVUJHZ89QkyL6cHvizZEB27AOLu
JqVZYiFMszcfkUAVYvs5SOxU5IRskNrS+YodN+2IeRjtJXesRSUszX30c2HAOHdMoXbDxllRJ3CO
NE42ollc3IopTd7mQqvWs376fknq7LJPrbqQrccPKeUbjUegbODcHslzroJB1BX90TpqiGW5UgYK
S1DSJlB2FRnhfJe+H5TFGGjWZaWEt8G0b4JSjfrrsVshMJEQYQV3Ap2yZSt/lxIpMHqdyVxyncwD
1Lwa4LNRvegt+3HwaQQu3LCtpdHxuqAJnoVV8dBt1hPYGWn94f2arAbIciH8dv9BY7ngJLstzvTv
eLI+IqZpN26i5+K46Tk4gwWLlT22nHRnxof455W4DAf2IQb1HXjKtXheF74FMXibFNgnRI4QfreR
0vA4lHu5zaxcRXYglVcrEvCtEyGYXUlTfQSZaE0aUBrpUhfOsv25InKDHjXWE2brm8FUlhRL3gBR
z/l6E4NV49jxW/t6JmWxemh2VN7oaRFMfR+Bgq5sdBV4Ndl4EfJoGXxej0zdmE1qV9drc6WsbZbP
w7SfQ7wCuequ131baXbZ7DLzvOnvfixFfGTkBcuieD2/vpXQFNzLOZe1wTCKGAufJLzp1sqxvShy
5P8Cg8i1AFSgynRonAAxDyV+sY5xyvmoI7k85j4NLHDea/s/Yxp8Misp4y7MkYK+nhSY7oAmD4mn
OuCfTdFs8apAyERAlUZtdwP5JXugojt4x0kEWFHTeSfDw9lMVmY8i9zyPsiKQrHvG7cffZdaPmmA
mYUmmxHXLLfA6EAi4nA+Ki9YXq2fHjjX8uBmjDurASLa114tPiVRXnwX4IJwDLpRT28h2JkU0lhg
tVI8RjDlhAkkyxrf7UpQuoygDfJIQnEX3mVSb81RJvVocxUaZMQUGWPEzYkBpcYoJ06e+hlugIIg
hRIROlVmJIik3G/xsG0jiZ8SMFimqELv+oGXgZ+V1WkNFk0RuleULdYf7362MM5z4EVP/aKcb7AX
fB8GzsdUE1bfZNuBbD5pbb22hnWulVzuloDa0RSjIEen3TR0yYm1h+CAk21pNckduIDP8BP4Cl9U
Ehg4fDROfW4WIGPNiEQza5opwrOY/FpH609Y3v95ol5JVxrYpWpsC20c7jh6ZgqvYndh/V/HPNf6
gE+m9H0xgzN95HF9lwshPbeaHgQP7E3pHApkGehP5bmrbz2ztpYxJdYUUlZJYxFpN833oq4UX4rE
GHvQcZxhqH48yN6MMu3q5m99yxDOEefVufjjXSnaxYyaS2e7pf8zG1dVUMPcbl6Iz1Wf+uMC05Fv
jaH9QLVy6410dtgk7o590EqX7WUMwfWiYZcVYAqsxDbp9FFjHxX5+3+5LN7p2lhpCKSQHAIPXGIo
SaylQNH/6/KOqiTZQu7d9vuD8W2MOt+PAOuCl4hHHm4dTz+L+JXx1594PWDp/fH8Yu720cvZrLV+
k9ybiPmMoAQCIeBGg0010AtzHmVQ0QSiKMN4vXg5gnDmMMhdWYciCsbARsHlvyEbv31UkXUKhAlZ
-- ==============================================================
-- RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
-- Version: 2020.1
-- Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
-- 
-- ===========================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity myproject is
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    fc1_input_V_ap_vld : IN STD_LOGIC;
    fc1_input_V : IN STD_LOGIC_VECTOR (111 downto 0);
    layer13_out_0_V : OUT STD_LOGIC_VECTOR (40 downto 0);
    layer13_out_0_V_ap_vld : OUT STD_LOGIC;
    layer13_out_1_V : OUT STD_LOGIC_VECTOR (40 downto 0);
    layer13_out_1_V_ap_vld : OUT STD_LOGIC;
    layer13_out_2_V : OUT STD_LOGIC_VECTOR (40 downto 0);
    layer13_out_2_V_ap_vld : OUT STD_LOGIC;
    layer13_out_3_V : OUT STD_LOGIC_VECTOR (40 downto 0);
    layer13_out_3_V_ap_vld : OUT STD_LOGIC;
    layer13_out_4_V : OUT STD_LOGIC_VECTOR (40 downto 0);
    layer13_out_4_V_ap_vld : OUT STD_LOGIC;
    const_size_in_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
    const_size_in_1_ap_vld : OUT STD_LOGIC;
    const_size_out_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
    const_size_out_1_ap_vld : OUT STD_LOGIC );
end;


architecture behav of myproject is 
    attribute CORE_GENERATION_INFO : STRING;
    attribute CORE_GENERATION_INFO of behav : architecture is
    "myproject,hls_ip_2020_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xcu250-figd2104-2L-e,HLS_INPUT_CLOCK=5.000000,HLS_INPUT_ARCH=pipeline,HLS_SYN_CLOCK=4.310000,HLS_SYN_LAT=10,HLS_SYN_TPT=1,HLS_SYN_MEM=4,HLS_SYN_DSP=5,HLS_SYN_FF=4312,HLS_SYN_LUT=47078,HLS_VERSION=2020_1}";
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';
    constant ap_ST_fsm_pp0_stage0 : STD_LOGIC_VECTOR (0 downto 0) := "1";
    constant ap_const_lv32_0 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000000";
    constant ap_const_boolean_1 : BOOLEAN := true;
    constant ap_const_boolean_0 : BOOLEAN := false;
    constant ap_const_lv112_0 : STD_LOGIC_VECTOR (111 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_const_lv16_10 : STD_LOGIC_VECTOR (15 downto 0) := "0000000000010000";
    constant ap_const_lv16_5 : STD_LOGIC_VECTOR (15 downto 0) := "0000000000000101";

    signal ap_CS_fsm : STD_LOGIC_VECTOR (0 downto 0) := "1";
    attribute fsm_encoding : string;
    attribute fsm_encoding of ap_CS_fsm : signal is "none";
    signal ap_CS_fsm_pp0_stage0 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage0 : signal is "none";
    signal ap_enable_reg_pp0_iter0 : STD_LOGIC;
    signal ap_enable_reg_pp0_iter1 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter2 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter3 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter4 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter5 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter6 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter7 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter8 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter9 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter10 : STD_LOGIC := '0';
    signal ap_idle_pp0 : STD_LOGIC;
    signal fc1_input_V_ap_vld_in_sig : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10 : BOOLEAN;
    signal ap_block_pp0_stage0_11001 : BOOLEAN;
    signal fc1_input_V_preg : STD_LOGIC_VECTOR (111 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    signal fc1_input_V_in_sig : STD_LOGIC_VECTOR (111 downto 0);
    signal fc1_input_V_ap_vld_preg : STD_LOGIC := '0';
    signal fc1_input_V_blk_n : STD_LOGIC;
    signal ap_block_pp0_stage0 : BOOLEAN;
    signal layer2_out_0_V_reg_1433 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_1_V_reg_1438 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_2_V_reg_1443 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_3_V_reg_1448 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_4_V_reg_1453 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_5_V_reg_1458 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_6_V_reg_1463 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_7_V_reg_1468 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_8_V_reg_1473 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_9_V_reg_1478 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_10_V_reg_1483 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_11_V_reg_1488 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_12_V_reg_1493 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_13_V_reg_1498 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_14_V_reg_1503 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_15_V_reg_1508 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_16_V_reg_1513 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_17_V_reg_1518 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_18_V_reg_1523 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_19_V_reg_1528 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_20_V_reg_1533 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_21_V_reg_1538 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_22_V_reg_1543 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_23_V_reg_1548 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_24_V_reg_1553 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_25_V_reg_1558 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_26_V_reg_1563 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_27_V_reg_1568 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_28_V_reg_1573 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_29_V_reg_1578 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_30_V_reg_1583 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_31_V_reg_1588 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_32_V_reg_1593 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_33_V_reg_1598 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_34_V_reg_1603 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_35_V_reg_1608 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_36_V_reg_1613 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_37_V_reg_1618 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_38_V_reg_1623 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_39_V_reg_1628 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_40_V_reg_1633 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_41_V_reg_1638 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_42_V_reg_1643 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_43_V_reg_1648 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_44_V_reg_1653 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_45_V_reg_1658 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_46_V_reg_1663 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_47_V_reg_1668 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_48_V_reg_1673 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_49_V_reg_1678 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_50_V_reg_1683 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_51_V_reg_1688 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_52_V_reg_1693 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_53_V_reg_1698 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_54_V_reg_1703 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_55_V_reg_1708 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_56_V_reg_1713 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_57_V_reg_1718 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_58_V_reg_1723 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_59_V_reg_1728 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_60_V_reg_1733 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_61_V_reg_1738 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_62_V_reg_1743 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_63_V_reg_1748 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_0_V_reg_1753 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_1_V_reg_1758 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_2_V_reg_1763 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_3_V_reg_1768 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_4_V_reg_1773 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_5_V_reg_1778 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_6_V_reg_1783 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_7_V_reg_1788 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_8_V_reg_1793 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_9_V_reg_1798 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_10_V_reg_1803 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_11_V_reg_1808 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_12_V_reg_1813 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_13_V_reg_1818 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_14_V_reg_1823 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_15_V_reg_1828 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_16_V_reg_1833 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_17_V_reg_1838 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_18_V_reg_1843 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_19_V_reg_1848 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_20_V_reg_1853 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_21_V_reg_1858 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_22_V_reg_1863 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_23_V_reg_1868 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_24_V_reg_1873 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_25_V_reg_1878 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_26_V_reg_1883 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_27_V_reg_1888 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_28_V_reg_1893 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_29_V_reg_1898 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_30_V_reg_1903 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_31_V_reg_1908 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_32_V_reg_1913 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_33_V_reg_1918 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_34_V_reg_1923 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_35_V_reg_1928 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_36_V_reg_1933 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_37_V_reg_1938 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_38_V_reg_1943 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_39_V_reg_1948 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_40_V_reg_1953 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_41_V_reg_1958 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_42_V_reg_1963 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_43_V_reg_1968 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_44_V_reg_1973 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_45_V_reg_1978 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_46_V_reg_1983 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_47_V_reg_1988 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_48_V_reg_1993 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_49_V_reg_1998 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_50_V_reg_2003 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_51_V_reg_2008 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_52_V_reg_2013 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_53_V_reg_2018 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_54_V_reg_2023 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_55_V_reg_2028 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_56_V_reg_2033 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_57_V_reg_2038 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_58_V_reg_2043 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_59_V_reg_2048 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_60_V_reg_2053 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_61_V_reg_2058 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_62_V_reg_2063 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_63_V_reg_2068 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_0_V_reg_2073 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_1_V_reg_2078 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_2_V_reg_2083 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_3_V_reg_2088 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_4_V_reg_2093 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_5_V_reg_2098 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_6_V_reg_2103 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_7_V_reg_2108 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_8_V_reg_2113 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_9_V_reg_2118 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_10_V_reg_2123 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_11_V_reg_2128 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_12_V_reg_2133 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_13_V_reg_2138 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_14_V_reg_2143 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_15_V_reg_2148 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_16_V_reg_2153 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_17_V_reg_2158 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_18_V_reg_2163 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_19_V_reg_2168 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_20_V_reg_2173 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_21_V_reg_2178 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_22_V_reg_2183 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_23_V_reg_2188 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_24_V_reg_2193 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_25_V_reg_2198 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_26_V_reg_2203 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_27_V_reg_2208 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_28_V_reg_2213 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_29_V_reg_2218 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_30_V_reg_2223 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_31_V_reg_2228 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer8_out_0_V_reg_2233 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_2_V_reg_2238 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_3_V_reg_2243 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_5_V_reg_2248 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_6_V_reg_2253 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_7_V_reg_2258 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_8_V_reg_2263 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_9_V_reg_2268 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_10_V_reg_2273 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_12_V_reg_2278 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_14_V_reg_2283 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_15_V_reg_2288 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_17_V_reg_2293 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_19_V_reg_2298 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_20_V_reg_2303 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_21_V_reg_2308 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_24_V_reg_2313 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_25_V_reg_2318 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_26_V_reg_2323 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_27_V_reg_2328 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_28_V_reg_2333 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_29_V_reg_2338 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_31_V_reg_2343 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_0_V_reg_2348 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_2_V_reg_2353 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_3_V_reg_2358 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_5_V_reg_2363 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_6_V_reg_2368 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_7_V_reg_2373 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_8_V_reg_2378 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_9_V_reg_2383 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_10_V_reg_2388 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_12_V_reg_2393 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_14_V_reg_2398 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_15_V_reg_2403 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_17_V_reg_2408 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_19_V_reg_2413 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_20_V_reg_2418 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_21_V_reg_2423 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_24_V_reg_2428 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_25_V_reg_2433 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_26_V_reg_2438 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_27_V_reg_2443 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_28_V_reg_2448 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_29_V_reg_2453 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer10_out_31_V_reg_2458 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer11_out_0_V_reg_2463 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer11_out_1_V_reg_2468 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer11_out_2_V_reg_2473 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer11_out_3_V_reg_2478 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer11_out_4_V_reg_2483 : STD_LOGIC_VECTOR (15 downto 0);
    signal ap_block_pp0_stage0_subdone : BOOLEAN;
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call145 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call145 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call145 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call145 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call145 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call145 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call145 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call145 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call145 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9_ignore_call145 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10_ignore_call145 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp143 : BOOLEAN;
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call211 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call211 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call211 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call211 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call211 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call211 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call211 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call211 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call211 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9_ignore_call211 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10_ignore_call211 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp210 : BOOLEAN;
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_ready : STD_LOGIC;
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_32 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_33 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_34 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_35 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_36 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_37 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_38 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_39 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_40 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_41 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_42 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_43 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_44 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_45 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_46 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_47 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_48 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_49 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_50 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_51 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_52 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_53 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_54 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_55 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_56 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_57 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_58 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_59 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_60 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_61 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_62 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_63 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_ready : STD_LOGIC;
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_0 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_1 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_2 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_3 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_4 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_5 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_6 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_7 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_8 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_9 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_10 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_11 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_12 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_13 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_14 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_15 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_16 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_17 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_18 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_19 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_20 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_21 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_22 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_23 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_24 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_25 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_26 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_27 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_28 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_29 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_30 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_31 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_32 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_33 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_34 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_35 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_36 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_37 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_38 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_39 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_40 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_41 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_42 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_43 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_44 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_45 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_46 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_47 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_48 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_49 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_50 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_51 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_52 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_53 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_54 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_55 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_56 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_57 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_58 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_59 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_60 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_61 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_62 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_63 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_ready : STD_LOGIC;
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_0 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_1 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_2 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_3 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_4 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_5 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_6 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_7 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_8 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_9 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_10 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_11 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_12 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_13 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_14 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_15 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_16 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_17 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_18 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_19 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_20 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_21 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_22 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_23 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_24 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_25 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_26 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_27 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_28 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_29 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_30 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_31 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_ready : STD_LOGIC;
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_0 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_1 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_2 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_3 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_4 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_5 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_6 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_7 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_8 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_9 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_10 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_11 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_12 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_13 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_14 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_15 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_16 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_17 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_18 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_19 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_20 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_21 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_22 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_ready : STD_LOGIC;
    signal call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_done : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_idle : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_ready : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_ce : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_0 : STD_LOGIC_VECTOR (40 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_1 : STD_LOGIC_VECTOR (40 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_2 : STD_LOGIC_VECTOR (40 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_3 : STD_LOGIC_VECTOR (40 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_4 : STD_LOGIC_VECTOR (40 downto 0);
    signal ap_block_state1_pp0_stage0_iter0_ignore_call265 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call265 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call265 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call265 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call265 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call265 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call265 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call265 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call265 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9_ignore_call265 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10_ignore_call265 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp265 : BOOLEAN;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start_reg : STD_LOGIC := '0';
    signal ap_block_pp0_stage0_01001 : BOOLEAN;
    signal ap_NS_fsm : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_idle_pp0_0to9 : STD_LOGIC;
    signal ap_reset_idle_pp0 : STD_LOGIC;
    signal ap_enable_pp0 : STD_LOGIC;

    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2 IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_32_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_33_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_34_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_35_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_36_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_37_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_38_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_39_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_40_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_41_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_42_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_43_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_44_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_45_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_46_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_47_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_48_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_49_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_50_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_51_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_52_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_53_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_54_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_55_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_56_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_57_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_58_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_59_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_60_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_61_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_62_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_63_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_V_read : IN STD_LOGIC_VECTOR (111 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_32 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_33 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_34 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_35 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_36 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_37 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_38 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_39 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_40 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_41 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_42 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_43 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_44 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_45 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_46 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_47 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_48 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_49 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_50 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_51 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_52 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_53 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_54 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_55 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_56 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_57 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_58 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_59 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_60 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_61 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_62 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_63 : OUT STD_LOGIC_VECTOR (15 downto 0) );
    end component;


    component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_32_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_33_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_34_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_35_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_36_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_37_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_38_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_39_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_40_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_41_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_42_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_43_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_44_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_45_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_46_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_47_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_48_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_49_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_50_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_51_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_52_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_53_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_54_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_55_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_56_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_57_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_58_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_59_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_60_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_61_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_62_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_63_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_32 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_33 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_34 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_35 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_36 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_37 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_38 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_39 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_40 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_41 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_42 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_43 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_44 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_45 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_46 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_47 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_48 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_49 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_50 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_51 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_52 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_53 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_54 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_55 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_56 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_57 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_58 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_59 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_60 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_61 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_62 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_63 : OUT STD_LOGIC_VECTOR (6 downto 0) );
    end component;


    component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (6 downto 0) );
    end component;


    component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (6 downto 0) );
    end component;


    component dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0 IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0) );
    end component;


    component softmax_latency_ap_fixed_ap_fixed_softmax_config13_s IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        ap_start : IN STD_LOGIC;
        ap_done : OUT STD_LOGIC;
        ap_idle : OUT STD_LOGIC;
        ap_ready : OUT STD_LOGIC;
        ap_ce : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (40 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (40 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (40 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (40 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (40 downto 0) );
    end component;



begin
    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_0_V_read => layer4_out_0_V_reg_1753,
        data_1_V_read => layer4_out_1_V_reg_1758,
        data_2_V_read => layer4_out_2_V_reg_1763,
        data_3_V_read => layer4_out_3_V_reg_1768,
        data_4_V_read => layer4_out_4_V_reg_1773,
        data_5_V_read => layer4_out_5_V_reg_1778,
        data_6_V_read => layer4_out_6_V_reg_1783,
        data_7_V_read => layer4_out_7_V_reg_1788,
        data_8_V_read => layer4_out_8_V_reg_1793,
        data_9_V_read => layer4_out_9_V_reg_1798,
        data_10_V_read => layer4_out_10_V_reg_1803,
        data_11_V_read => layer4_out_11_V_reg_1808,
        data_12_V_read => layer4_out_12_V_reg_1813,
        data_13_V_read => layer4_out_13_V_reg_1818,
        data_14_V_read => layer4_out_14_V_reg_1823,
        data_15_V_read => layer4_out_15_V_reg_1828,
        data_16_V_read => layer4_out_16_V_reg_1833,
        data_17_V_read => layer4_out_17_V_reg_1838,
        data_18_V_read => layer4_out_18_V_reg_1843,
        data_19_V_read => layer4_out_19_V_reg_1848,
        data_20_V_read => layer4_out_20_V_reg_1853,
        data_21_V_read => layer4_out_21_V_reg_1858,
        data_22_V_read => layer4_out_22_V_reg_1863,
        data_23_V_read => layer4_out_23_V_reg_1868,
        data_24_V_read => layer4_out_24_V_reg_1873,
        data_25_V_read => layer4_out_25_V_reg_1878,
        data_26_V_read => layer4_out_26_V_reg_1883,
        data_27_V_read => layer4_out_27_V_reg_1888,
        data_28_V_read => layer4_out_28_V_reg_1893,
        data_29_V_read => layer4_out_29_V_reg_1898,
        data_30_V_read => layer4_out_30_V_reg_1903,
        data_31_V_read => layer4_out_31_V_reg_1908,
        data_32_V_read => layer4_out_32_V_reg_1913,
        data_33_V_read => layer4_out_33_V_reg_1918,
        data_34_V_read => layer4_out_34_V_reg_1923,
        data_35_V_read => layer4_out_35_V_reg_1928,
        data_36_V_read => layer4_out_36_V_reg_1933,
        data_37_V_read => layer4_out_37_V_reg_1938,
        data_38_V_read => layer4_out_38_V_reg_1943,
        data_39_V_read => layer4_out_39_V_reg_1948,
        data_40_V_read => layer4_out_40_V_reg_1953,
        data_41_V_read => layer4_out_41_V_reg_1958,
        data_42_V_read => layer4_out_42_V_reg_1963,
        data_43_V_read => layer4_out_43_V_reg_1968,
        data_44_V_read => layer4_out_44_V_reg_1973,
        data_45_V_read => layer4_out_45_V_reg_1978,
        data_46_V_read => layer4_out_46_V_reg_1983,
        data_47_V_read => layer4_out_47_V_reg_1988,
        data_48_V_read => layer4_out_48_V_reg_1993,
        data_49_V_read => layer4_out_49_V_reg_1998,
        data_50_V_read => layer4_out_50_V_reg_2003,
        data_51_V_read => layer4_out_51_V_reg_2008,
        data_52_V_read => layer4_out_52_V_reg_2013,
        data_53_V_read => layer4_out_53_V_reg_2018,
        data_54_V_read => layer4_out_54_V_reg_2023,
        data_55_V_read => layer4_out_55_V_reg_2028,
        data_56_V_read => layer4_out_56_V_reg_2033,
        data_57_V_read => layer4_out_57_V_reg_2038,
        data_58_V_read => layer4_out_58_V_reg_2043,
        data_59_V_read => layer4_out_59_V_reg_2048,
        data_60_V_read => layer4_out_60_V_reg_2053,
        data_61_V_read => layer4_out_61_V_reg_2058,
        data_62_V_read => layer4_out_62_V_reg_2063,
        data_63_V_read => layer4_out_63_V_reg_2068,
        ap_return_0 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_0,
        ap_return_1 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_1,
        ap_return_2 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_2,
        ap_return_3 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_3,
        ap_return_4 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_4,
        ap_return_5 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_5,
        ap_return_6 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_6,
        ap_return_7 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_7,
        ap_return_8 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_8,
        ap_return_9 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_9,
        ap_return_10 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_10,
        ap_return_11 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_11,
        ap_return_12 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_12,
        ap_return_13 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_13,
        ap_return_14 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_14,
        ap_return_15 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_15,
        ap_return_16 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_16,
        ap_return_17 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_17,
        ap_return_18 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_18,
        ap_return_19 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_19,
        ap_return_20 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_20,
        ap_return_21 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_21,
        ap_return_22 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_22,
        ap_return_23 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_23,
        ap_return_24 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_24,
        ap_return_25 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_25,
        ap_return_26 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_26,
        ap_return_27 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_27,
        ap_return_28 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_28,
        ap_return_29 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_29,
        ap_return_30 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_30,
        ap_return_31 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_31,
        ap_ce => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_ce);

    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_0_V_read => layer7_out_0_V_reg_2073,
        data_1_V_read => layer7_out_1_V_reg_2078,
        data_2_V_read => layer7_out_2_V_reg_2083,
        data_3_V_read => layer7_out_3_V_reg_2088,
        data_4_V_read => layer7_out_4_V_reg_2093,
        data_5_V_read => layer7_out_5_V_reg_2098,
        data_6_V_read => layer7_out_6_V_reg_2103,
        data_7_V_read => layer7_out_7_V_reg_2108,
        data_8_V_read => layer7_out_8_V_reg_2113,
        data_9_V_read => layer7_out_9_V_reg_2118,
        data_10_V_read => layer7_out_10_V_reg_2123,
        data_11_V_read => layer7_out_11_V_reg_2128,
        data_12_V_read => layer7_out_12_V_reg_2133,
        data_13_V_read => layer7_out_13_V_reg_2138,
        data_14_V_read => layer7_out_14_V_reg_2143,
        data_15_V_read => layer7_out_15_V_reg_2148,
        data_16_V_read => layer7_out_16_V_reg_2153,
        data_17_V_read => layer7_out_17_V_reg_2158,
        data_18_V_read => layer7_out_18_V_reg_2163,
        data_19_V_read => layer7_out_19_V_reg_2168,
        data_20_V_read => layer7_out_20_V_reg_2173,
        data_21_V_read => layer7_out_21_V_reg_2178,
        data_22_V_read => layer7_out_22_V_reg_2183,
        data_23_V_read => layer7_out_23_V_reg_2188,
        data_24_V_read => layer7_out_24_V_reg_2193,
        data_25_V_read => layer7_out_25_V_reg_2198,
        data_26_V_read => layer7_out_26_V_reg_2203,
        data_27_V_read => layer7_out_27_V_reg_2208,
        data_28_V_read => layer7_out_28_V_reg_2213,
        data_29_V_read => layer7_out_29_V_reg_2218,
        data_30_V_read => layer7_out_30_V_reg_2223,
        data_31_V_read => layer7_out_31_V_reg_2228,
        ap_return_0 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_0,
        ap_return_1 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_1,
        ap_return_2 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_2,
        ap_return_3 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_3,
        ap_return_4 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_4,
        ap_return_5 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_5,
        ap_return_6 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_6,
        ap_return_7 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_7,
        ap_return_8 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_8,
        ap_return_9 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_9,
        ap_return_10 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_10,
        ap_return_11 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_11,
        ap_return_12 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_12,
        ap_return_13 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_13,
        ap_return_14 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_14,
        ap_return_15 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_15,
        ap_return_16 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_16,
        ap_return_17 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_17,
        ap_return_18 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_18,
        ap_return_19 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_19,
        ap_return_20 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_20,
        ap_return_21 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_21,
        ap_return_22 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_22,
        ap_ce => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_ce);

    call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s
    port map (
        ap_ready => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_ready,
        data_V_read => fc1_input_V_in_sig,
        ap_return_0 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_0,
        ap_return_1 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_1,
        ap_return_2 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_2,
        ap_return_3 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_3,
        ap_return_4 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_4,
        ap_return_5 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_5,
        ap_return_6 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_6,
        ap_return_7 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_7,
        ap_return_8 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_8,
        ap_return_9 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_9,
        ap_return_10 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_10,
        ap_return_11 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_11,
        ap_return_12 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_12,
        ap_return_13 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_13,
        ap_return_14 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_14,
        ap_return_15 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_15,
        ap_return_16 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_16,
        ap_return_17 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_17,
        ap_return_18 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_18,
        ap_return_19 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_19,
        ap_return_20 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_20,
        ap_return_21 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_21,
        ap_return_22 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_22,
        ap_return_23 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_23,
        ap_return_24 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_24,
        ap_return_25 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_25,
        ap_return_26 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_26,
        ap_return_27 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_27,
        ap_return_28 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_28,
        ap_return_29 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_29,
        ap_return_30 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_30,
        ap_return_31 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_31,
        ap_return_32 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_32,
        ap_return_33 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_33,
        ap_return_34 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_34,
        ap_return_35 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_35,
        ap_return_36 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_36,
        ap_return_37 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_37,
        ap_return_38 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_38,
        ap_return_39 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_39,
        ap_return_40 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_40,
        ap_return_41 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_41,
        ap_return_42 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_42,
        ap_return_43 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_43,
        ap_return_44 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_44,
        ap_return_45 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_45,
        ap_return_46 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_46,
        ap_return_47 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_47,
        ap_return_48 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_48,
        ap_return_49 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_49,
        ap_return_50 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_50,
        ap_return_51 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_51,
        ap_return_52 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_52,
        ap_return_53 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_53,
        ap_return_54 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_54,
        ap_return_55 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_55,
        ap_return_56 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_56,
        ap_return_57 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_57,
        ap_return_58 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_58,
        ap_return_59 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_59,
        ap_return_60 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_60,
        ap_return_61 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_61,
        ap_return_62 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_62,
        ap_return_63 => call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_63);

    call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233 : component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s
    port map (
        ap_ready => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_ready,
        data_0_V_read => layer2_out_0_V_reg_1433,
        data_1_V_read => layer2_out_1_V_reg_1438,
        data_2_V_read => layer2_out_2_V_reg_1443,
        data_3_V_read => layer2_out_3_V_reg_1448,
        data_4_V_read => layer2_out_4_V_reg_1453,
        data_5_V_read => layer2_out_5_V_reg_1458,
        data_6_V_read => layer2_out_6_V_reg_1463,
        data_7_V_read => layer2_out_7_V_reg_1468,
        data_8_V_read => layer2_out_8_V_reg_1473,
        data_9_V_read => layer2_out_9_V_reg_1478,
        data_10_V_read => layer2_out_10_V_reg_1483,
        data_11_V_read => layer2_out_11_V_reg_1488,
        data_12_V_read => layer2_out_12_V_reg_1493,
        data_13_V_read => layer2_out_13_V_reg_1498,
        data_14_V_read => layer2_out_14_V_reg_1503,
        data_15_V_read => layer2_out_15_V_reg_1508,
        data_16_V_read => layer2_out_16_V_reg_1513,
        data_17_V_read => layer2_out_17_V_reg_1518,
        data_18_V_read => layer2_out_18_V_reg_1523,
        data_19_V_read => layer2_out_19_V_reg_1528,
        data_20_V_read => layer2_out_20_V_reg_1533,
        data_21_V_read => layer2_out_21_V_reg_1538,
        data_22_V_read => layer2_out_22_V_reg_1543,
        data_23_V_read => layer2_out_23_V_reg_1548,
        data_24_V_read => layer2_out_24_V_reg_1553,
        data_25_V_read => layer2_out_25_V_reg_1558,
        data_26_V_read => layer2_out_26_V_reg_1563,
        data_27_V_read => layer2_out_27_V_reg_1568,
        data_28_V_read => layer2_out_28_V_reg_1573,
        data_29_V_read => layer2_out_29_V_reg_1578,
        data_30_V_read => layer2_out_30_V_reg_1583,
        data_31_V_read => layer2_out_31_V_reg_1588,
        data_32_V_read => layer2_out_32_V_reg_1593,
        data_33_V_read => layer2_out_33_V_reg_1598,
        data_34_V_read => layer2_out_34_V_reg_1603,
        data_35_V_read => layer2_out_35_V_reg_1608,
        data_36_V_read => layer2_out_36_V_reg_1613,
        data_37_V_read => layer2_out_37_V_reg_1618,
        data_38_V_read => layer2_out_38_V_reg_1623,
        data_39_V_read => layer2_out_39_V_reg_1628,
        data_40_V_read => layer2_out_40_V_reg_1633,
        data_41_V_read => layer2_out_41_V_reg_1638,
        data_42_V_read => layer2_out_42_V_reg_1643,
        data_43_V_read => layer2_out_43_V_reg_1648,
        data_44_V_read => layer2_out_44_V_reg_1653,
        data_45_V_read => layer2_out_45_V_reg_1658,
        data_46_V_read => layer2_out_46_V_reg_1663,
        data_47_V_read => layer2_out_47_V_reg_1668,
        data_48_V_read => layer2_out_48_V_reg_1673,
        data_49_V_read => layer2_out_49_V_reg_1678,
        data_50_V_read => layer2_out_50_V_reg_1683,
        data_51_V_read => layer2_out_51_V_reg_1688,
        data_52_V_read => layer2_out_52_V_reg_1693,
        data_53_V_read => layer2_out_53_V_reg_1698,
        data_54_V_read => layer2_out_54_V_reg_1703,
        data_55_V_read => layer2_out_55_V_reg_1708,
        data_56_V_read => layer2_out_56_V_reg_1713,
        data_57_V_read => layer2_out_57_V_reg_1718,
        data_58_V_read => layer2_out_58_V_reg_1723,
        data_59_V_read => layer2_out_59_V_reg_1728,
        data_60_V_read => layer2_out_60_V_reg_1733,
        data_61_V_read => layer2_out_61_V_reg_1738,
        data_62_V_read => layer2_out_62_V_reg_1743,
        data_63_V_read => layer2_out_63_V_reg_1748,
        ap_return_0 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_0,
        ap_return_1 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_1,
        ap_return_2 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_2,
        ap_return_3 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_3,
        ap_return_4 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_4,
        ap_return_5 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_5,
        ap_return_6 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_6,
        ap_return_7 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_7,
        ap_return_8 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_8,
        ap_return_9 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_9,
        ap_return_10 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_10,
        ap_return_11 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_11,
        ap_return_12 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_12,
        ap_return_13 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_13,
        ap_return_14 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_14,
        ap_return_15 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_15,
        ap_return_16 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_16,
        ap_return_17 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_17,
        ap_return_18 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_18,
        ap_return_19 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_19,
        ap_return_20 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_20,
        ap_return_21 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_21,
        ap_return_22 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_22,
        ap_return_23 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_23,
        ap_return_24 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_24,
        ap_return_25 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_25,
        ap_return_26 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_26,
        ap_return_27 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_27,
        ap_return_28 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_28,
        ap_return_29 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_29,
        ap_return_30 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_30,
        ap_return_31 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_31,
        ap_return_32 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_32,
        ap_return_33 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_33,
        ap_return_34 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_34,
        ap_return_35 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_35,
        ap_return_36 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_36,
        ap_return_37 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_37,
        ap_return_38 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_38,
        ap_return_39 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_39,
        ap_return_40 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_40,
        ap_return_41 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_41,
        ap_return_42 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_42,
        ap_return_43 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_43,
        ap_return_44 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_44,
        ap_return_45 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_45,
        ap_return_46 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_46,
        ap_return_47 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_47,
        ap_return_48 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_48,
        ap_return_49 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_49,
        ap_return_50 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_50,
        ap_return_51 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_51,
        ap_return_52 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_52,
        ap_return_53 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_53,
        ap_return_54 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_54,
        ap_return_55 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_55,
        ap_return_56 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_56,
        ap_return_57 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_57,
        ap_return_58 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_58,
        ap_return_59 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_59,
        ap_return_60 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_60,
        ap_return_61 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_61,
        ap_return_62 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_62,
        ap_return_63 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_63);

    call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301 : component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s
    port map (
        ap_ready => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_ready,
        data_0_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_0,
        data_1_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_1,
        data_2_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_2,
        data_3_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_3,
        data_4_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_4,
        data_5_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_5,
        data_6_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_6,
        data_7_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_7,
        data_8_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_8,
        data_9_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_9,
        data_10_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_10,
        data_11_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_11,
        data_12_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_12,
        data_13_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_13,
        data_14_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_14,
        data_15_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_15,
        data_16_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_16,
        data_17_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_17,
        data_18_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_18,
        data_19_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_19,
        data_20_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_20,
        data_21_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_21,
        data_22_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_22,
        data_23_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_23,
        data_24_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_24,
        data_25_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_25,
        data_26_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_26,
        data_27_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_27,
        data_28_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_28,
        data_29_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_29,
        data_30_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_30,
        data_31_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_return_31,
        ap_return_0 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_0,
        ap_return_1 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_1,
        ap_return_2 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_2,
        ap_return_3 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_3,
        ap_return_4 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_4,
        ap_return_5 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_5,
        ap_return_6 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_6,
        ap_return_7 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_7,
        ap_return_8 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_8,
        ap_return_9 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_9,
        ap_return_10 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_10,
        ap_return_11 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_11,
        ap_return_12 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_12,
        ap_return_13 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_13,
        ap_return_14 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_14,
        ap_return_15 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_15,
        ap_return_16 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_16,
        ap_return_17 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_17,
        ap_return_18 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_18,
        ap_return_19 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_19,
        ap_return_20 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_20,
        ap_return_21 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_21,
        ap_return_22 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_22,
        ap_return_23 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_23,
        ap_return_24 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_24,
        ap_return_25 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_25,
        ap_return_26 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_26,
        ap_return_27 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_27,
        ap_return_28 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_28,
        ap_return_29 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_29,
        ap_return_30 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_30,
        ap_return_31 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_31);

    call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337 : component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s
    port map (
        ap_ready => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_ready,
        data_0_V_read => layer8_out_0_V_reg_2233,
        data_2_V_read => layer8_out_2_V_reg_2238,
        data_3_V_read => layer8_out_3_V_reg_2243,
        data_5_V_read => layer8_out_5_V_reg_2248,
        data_6_V_read => layer8_out_6_V_reg_2253,
        data_7_V_read => layer8_out_7_V_reg_2258,
        data_8_V_read => layer8_out_8_V_reg_2263,
        data_9_V_read => layer8_out_9_V_reg_2268,
        data_10_V_read => layer8_out_10_V_reg_2273,
        data_12_V_read => layer8_out_12_V_reg_2278,
        data_14_V_read => layer8_out_14_V_reg_2283,
        data_15_V_read => layer8_out_15_V_reg_2288,
        data_17_V_read => layer8_out_17_V_reg_2293,
        data_19_V_read => layer8_out_19_V_reg_2298,
        data_20_V_read => layer8_out_20_V_reg_2303,
        data_21_V_read => layer8_out_21_V_reg_2308,
        data_24_V_read => layer8_out_24_V_reg_2313,
        data_25_V_read => layer8_out_25_V_reg_2318,
        data_26_V_read => layer8_out_26_V_reg_2323,
        data_27_V_read => layer8_out_27_V_reg_2328,
        data_28_V_read => layer8_out_28_V_reg_2333,
        data_29_V_read => layer8_out_29_V_reg_2338,
        data_31_V_read => layer8_out_31_V_reg_2343,
        ap_return_0 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_0,
        ap_return_1 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_1,
        ap_return_2 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_2,
        ap_return_3 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_3,
        ap_return_4 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_4,
        ap_return_5 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_5,
        ap_return_6 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_6,
        ap_return_7 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_7,
        ap_return_8 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_8,
        ap_return_9 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_9,
        ap_return_10 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_10,
        ap_return_11 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_11,
        ap_return_12 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_12,
        ap_return_13 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_13,
        ap_return_14 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_14,
        ap_return_15 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_15,
        ap_return_16 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_16,
        ap_return_17 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_17,
        ap_return_18 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_18,
        ap_return_19 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_19,
        ap_return_20 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_20,
        ap_return_21 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_21,
        ap_return_22 => call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_22);

    call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364 : component dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0
    port map (
        ap_ready => call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_ready,
        data_0_V_read => layer10_out_0_V_reg_2348,
        data_2_V_read => layer10_out_2_V_reg_2353,
        data_3_V_read => layer10_out_3_V_reg_2358,
        data_5_V_read => layer10_out_5_V_reg_2363,
        data_6_V_read => layer10_out_6_V_reg_2368,
        data_7_V_read => layer10_out_7_V_reg_2373,
        data_8_V_read => layer10_out_8_V_reg_2378,
        data_9_V_read => layer10_out_9_V_reg_2383,
        data_10_V_read => layer10_out_10_V_reg_2388,
        data_12_V_read => layer10_out_12_V_reg_2393,
        data_14_V_read => layer10_out_14_V_reg_2398,
        data_15_V_read => layer10_out_15_V_reg_2403,
        data_17_V_read => layer10_out_17_V_reg_2408,
        data_19_V_read => layer10_out_19_V_reg_2413,
        data_20_V_read => layer10_out_20_V_reg_2418,
        data_21_V_read => layer10_out_21_V_reg_2423,
        data_24_V_read => layer10_out_24_V_reg_2428,
        data_25_V_read => layer10_out_25_V_reg_2433,
        data_26_V_read => layer10_out_26_V_reg_2438,
        data_27_V_read => layer10_out_27_V_reg_2443,
        data_28_V_read => layer10_out_28_V_reg_2448,
        data_29_V_read => layer10_out_29_V_reg_2453,
        data_31_V_read => layer10_out_31_V_reg_2458,
        ap_return_0 => call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_0,
        ap_return_1 => call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_1,
        ap_return_2 => call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_2,
        ap_return_3 => call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_3,
        ap_return_4 => call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_4);

    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391 : component softmax_latency_ap_fixed_ap_fixed_softmax_config13_s
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        ap_start => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start,
        ap_done => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_done,
        ap_idle => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_idle,
        ap_ready => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_ready,
        ap_ce => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_ce,
        data_0_V_read => layer11_out_0_V_reg_2463,
        data_1_V_read => layer11_out_1_V_reg_2468,
        data_2_V_read => layer11_out_2_V_reg_2473,
        data_3_V_read => layer11_out_3_V_reg_2478,
        data_4_V_read => layer11_out_4_V_reg_2483,
        ap_return_0 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_0,
        ap_return_1 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_1,
        ap_return_2 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_2,
        ap_return_3 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_3,
        ap_return_4 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_4);





    ap_CS_fsm_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
            else
                ap_CS_fsm <= ap_NS_fsm;
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter1_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter1 <= ap_const_logic_0;
            else
                if (((ap_const_boolean_0 = ap_block_pp0_stage0_subdone) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
                    ap_enable_reg_pp0_iter1 <= ap_start;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter10_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter10 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter2_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter2 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter3_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter3 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter4_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter4 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter5_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter5 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter6_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter6 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter7_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter7 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter8_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter8 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter9_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter9 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
                end if; 
            end if;
        end if;
    end process;


    fc1_input_V_ap_vld_preg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                fc1_input_V_ap_vld_preg <= ap_const_logic_0;
            else
                if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
                    fc1_input_V_ap_vld_preg <= ap_const_logic_0;
                elsif ((not(((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) and (fc1_input_V_ap_vld = ap_const_logic_1))) then 
                    fc1_input_V_ap_vld_preg <= fc1_input_V_ap_vld;
                end if; 
            end if;
        end if;
    end process;


    fc1_input_V_preg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                fc1_input_V_preg <= ap_const_lv112_0;
            else
                if ((not(((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) and (fc1_input_V_ap_vld = ap_const_logic_1))) then 
                    fc1_input_V_preg <= fc1_input_V;
                end if; 
            end if;
        end if;
    end process;


    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start_reg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start_reg <= ap_const_logic_0;
            else
                if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter7 = ap_const_logic_1))) then 
                    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start_reg <= ap_const_logic_1;
                elsif ((grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_ready = ap_const_logic_1)) then 
                    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start_reg <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;

    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_const_boolean_0 = ap_block_pp0_stage0_11001)) then
                layer10_out_0_V_reg_2348 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_0;
                layer10_out_10_V_reg_2388 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_8;
                layer10_out_12_V_reg_2393 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_9;
                layer10_out_14_V_reg_2398 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_10;
                layer10_out_15_V_reg_2403 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_11;
                layer10_out_17_V_reg_2408 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_12;
                layer10_out_19_V_reg_2413 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_13;
                layer10_out_20_V_reg_2418 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_14;
                layer10_out_21_V_reg_2423 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_15;
                layer10_out_24_V_reg_2428 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_16;
                layer10_out_25_V_reg_2433 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_17;
                layer10_out_26_V_reg_2438 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_18;
                layer10_out_27_V_reg_2443 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_19;
                layer10_out_28_V_reg_2448 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_20;
                layer10_out_29_V_reg_2453 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_21;
                layer10_out_2_V_reg_2353 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_1;
                layer10_out_31_V_reg_2458 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_22;
                layer10_out_3_V_reg_2358 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_2;
                layer10_out_5_V_reg_2363 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_3;
                layer10_out_6_V_reg_2368 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_4;
                layer10_out_7_V_reg_2373 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_5;
                layer10_out_8_V_reg_2378 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_6;
                layer10_out_9_V_reg_2383 <= call_ret5_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config10_s_fu_337_ap_return_7;
                layer11_out_0_V_reg_2463 <= call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_0;
                layer11_out_1_V_reg_2468 <= call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_1;
                layer11_out_2_V_reg_2473 <= call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_2;
                layer11_out_3_V_reg_2478 <= call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_3;
                layer11_out_4_V_reg_2483 <= call_ret6_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_364_ap_return_4;
                layer7_out_0_V_reg_2073 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_0;
                layer7_out_10_V_reg_2123 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_10;
                layer7_out_11_V_reg_2128 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_11;
                layer7_out_12_V_reg_2133 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_12;
                layer7_out_13_V_reg_2138 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_13;
                layer7_out_14_V_reg_2143 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_14;
                layer7_out_15_V_reg_2148 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_15;
                layer7_out_16_V_reg_2153 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_16;
                layer7_out_17_V_reg_2158 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_17;
                layer7_out_18_V_reg_2163 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_18;
                layer7_out_19_V_reg_2168 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_19;
                layer7_out_1_V_reg_2078 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_1;
                layer7_out_20_V_reg_2173 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_20;
                layer7_out_21_V_reg_2178 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_21;
                layer7_out_22_V_reg_2183 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_22;
                layer7_out_23_V_reg_2188 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_23;
                layer7_out_24_V_reg_2193 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_24;
                layer7_out_25_V_reg_2198 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_25;
                layer7_out_26_V_reg_2203 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_26;
                layer7_out_27_V_reg_2208 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_27;
                layer7_out_28_V_reg_2213 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_28;
                layer7_out_29_V_reg_2218 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_29;
                layer7_out_2_V_reg_2083 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_2;
                layer7_out_30_V_reg_2223 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_30;
                layer7_out_31_V_reg_2228 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_31;
                layer7_out_3_V_reg_2088 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_3;
                layer7_out_4_V_reg_2093 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_4;
                layer7_out_5_V_reg_2098 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_5;
                layer7_out_6_V_reg_2103 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_6;
                layer7_out_7_V_reg_2108 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_7;
                layer7_out_8_V_reg_2113 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_8;
                layer7_out_9_V_reg_2118 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_301_ap_return_9;
                layer8_out_0_V_reg_2233 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_0;
                layer8_out_10_V_reg_2273 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_8;
                layer8_out_12_V_reg_2278 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_9;
                layer8_out_14_V_reg_2283 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_10;
                layer8_out_15_V_reg_2288 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_11;
                layer8_out_17_V_reg_2293 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_12;
                layer8_out_19_V_reg_2298 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_13;
                layer8_out_20_V_reg_2303 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_14;
                layer8_out_21_V_reg_2308 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_15;
                layer8_out_24_V_reg_2313 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_16;
                layer8_out_25_V_reg_2318 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_17;
                layer8_out_26_V_reg_2323 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_18;
                layer8_out_27_V_reg_2328 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_19;
                layer8_out_28_V_reg_2333 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_20;
                layer8_out_29_V_reg_2338 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_21;
                layer8_out_2_V_reg_2238 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_1;
                layer8_out_31_V_reg_2343 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_22;
                layer8_out_3_V_reg_2243 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_2;
                layer8_out_5_V_reg_2248 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_3;
                layer8_out_6_V_reg_2253 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_4;
                layer8_out_7_V_reg_2258 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_5;
                layer8_out_8_V_reg_2263 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_6;
                layer8_out_9_V_reg_2268 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_return_7;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then
                layer2_out_0_V_reg_1433 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_0;
                layer2_out_10_V_reg_1483 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_10;
                layer2_out_11_V_reg_1488 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_11;
                layer2_out_12_V_reg_1493 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_12;
                layer2_out_13_V_reg_1498 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_13;
                layer2_out_14_V_reg_1503 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_14;
                layer2_out_15_V_reg_1508 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_15;
                layer2_out_16_V_reg_1513 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_16;
                layer2_out_17_V_reg_1518 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_17;
                layer2_out_18_V_reg_1523 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_18;
                layer2_out_19_V_reg_1528 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_19;
                layer2_out_1_V_reg_1438 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_1;
                layer2_out_20_V_reg_1533 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_20;
                layer2_out_21_V_reg_1538 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_21;
                layer2_out_22_V_reg_1543 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_22;
                layer2_out_23_V_reg_1548 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_23;
                layer2_out_24_V_reg_1553 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_24;
                layer2_out_25_V_reg_1558 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_25;
                layer2_out_26_V_reg_1563 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_26;
                layer2_out_27_V_reg_1568 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_27;
                layer2_out_28_V_reg_1573 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_28;
                layer2_out_29_V_reg_1578 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_29;
                layer2_out_2_V_reg_1443 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_2;
                layer2_out_30_V_reg_1583 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_30;
                layer2_out_31_V_reg_1588 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_31;
                layer2_out_32_V_reg_1593 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_32;
                layer2_out_33_V_reg_1598 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_33;
                layer2_out_34_V_reg_1603 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_34;
                layer2_out_35_V_reg_1608 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_35;
                layer2_out_36_V_reg_1613 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_36;
                layer2_out_37_V_reg_1618 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_37;
                layer2_out_38_V_reg_1623 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_38;
                layer2_out_39_V_reg_1628 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_39;
                layer2_out_3_V_reg_1448 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_3;
                layer2_out_40_V_reg_1633 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_40;
                layer2_out_41_V_reg_1638 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_41;
                layer2_out_42_V_reg_1643 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_42;
                layer2_out_43_V_reg_1648 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_43;
                layer2_out_44_V_reg_1653 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_44;
                layer2_out_45_V_reg_1658 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_45;
                layer2_out_46_V_reg_1663 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_46;
                layer2_out_47_V_reg_1668 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_47;
                layer2_out_48_V_reg_1673 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_48;
                layer2_out_49_V_reg_1678 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_49;
                layer2_out_4_V_reg_1453 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_4;
                layer2_out_50_V_reg_1683 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_50;
                layer2_out_51_V_reg_1688 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_51;
                layer2_out_52_V_reg_1693 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_52;
                layer2_out_53_V_reg_1698 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_53;
                layer2_out_54_V_reg_1703 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_54;
                layer2_out_55_V_reg_1708 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_55;
                layer2_out_56_V_reg_1713 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_56;
                layer2_out_57_V_reg_1718 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_57;
                layer2_out_58_V_reg_1723 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_58;
                layer2_out_59_V_reg_1728 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_59;
                layer2_out_5_V_reg_1458 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_5;
                layer2_out_60_V_reg_1733 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_60;
                layer2_out_61_V_reg_1738 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_61;
                layer2_out_62_V_reg_1743 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_62;
                layer2_out_63_V_reg_1748 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_63;
                layer2_out_6_V_reg_1463 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_6;
                layer2_out_7_V_reg_1468 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_7;
                layer2_out_8_V_reg_1473 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_8;
                layer2_out_9_V_reg_1478 <= call_ret_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_227_ap_return_9;
                layer4_out_0_V_reg_1753 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_0;
                layer4_out_10_V_reg_1803 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_10;
                layer4_out_11_V_reg_1808 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_11;
                layer4_out_12_V_reg_1813 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_12;
                layer4_out_13_V_reg_1818 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_13;
                layer4_out_14_V_reg_1823 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_14;
                layer4_out_15_V_reg_1828 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_15;
                layer4_out_16_V_reg_1833 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_16;
                layer4_out_17_V_reg_1838 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_17;
                layer4_out_18_V_reg_1843 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_18;
                layer4_out_19_V_reg_1848 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_19;
                layer4_out_1_V_reg_1758 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_1;
                layer4_out_20_V_reg_1853 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_20;
                layer4_out_21_V_reg_1858 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_21;
                layer4_out_22_V_reg_1863 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_22;
                layer4_out_23_V_reg_1868 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_23;
                layer4_out_24_V_reg_1873 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_24;
                layer4_out_25_V_reg_1878 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_25;
                layer4_out_26_V_reg_1883 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_26;
                layer4_out_27_V_reg_1888 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_27;
                layer4_out_28_V_reg_1893 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_28;
                layer4_out_29_V_reg_1898 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_29;
                layer4_out_2_V_reg_1763 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_2;
                layer4_out_30_V_reg_1903 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_30;
                layer4_out_31_V_reg_1908 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_31;
                layer4_out_32_V_reg_1913 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_32;
                layer4_out_33_V_reg_1918 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_33;
                layer4_out_34_V_reg_1923 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_34;
                layer4_out_35_V_reg_1928 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_35;
                layer4_out_36_V_reg_1933 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_36;
                layer4_out_37_V_reg_1938 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_37;
                layer4_out_38_V_reg_1943 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_38;
                layer4_out_39_V_reg_1948 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_39;
                layer4_out_3_V_reg_1768 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_3;
                layer4_out_40_V_reg_1953 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_40;
                layer4_out_41_V_reg_1958 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_41;
                layer4_out_42_V_reg_1963 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_42;
                layer4_out_43_V_reg_1968 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_43;
                layer4_out_44_V_reg_1973 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_44;
                layer4_out_45_V_reg_1978 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_45;
                layer4_out_46_V_reg_1983 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_46;
                layer4_out_47_V_reg_1988 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_47;
                layer4_out_48_V_reg_1993 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_48;
                layer4_out_49_V_reg_1998 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_49;
                layer4_out_4_V_reg_1773 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_4;
                layer4_out_50_V_reg_2003 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_50;
                layer4_out_51_V_reg_2008 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_51;
                layer4_out_52_V_reg_2013 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_52;
                layer4_out_53_V_reg_2018 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_53;
                layer4_out_54_V_reg_2023 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_54;
                layer4_out_55_V_reg_2028 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_55;
                layer4_out_56_V_reg_2033 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_56;
                layer4_out_57_V_reg_2038 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_57;
                layer4_out_58_V_reg_2043 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_58;
                layer4_out_59_V_reg_2048 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_59;
                layer4_out_5_V_reg_1778 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_5;
                layer4_out_60_V_reg_2053 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_60;
                layer4_out_61_V_reg_2058 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_61;
                layer4_out_62_V_reg_2063 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_62;
                layer4_out_63_V_reg_2068 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_63;
                layer4_out_6_V_reg_1783 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_6;
                layer4_out_7_V_reg_1788 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_7;
                layer4_out_8_V_reg_1793 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_8;
                layer4_out_9_V_reg_1798 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_233_ap_return_9;
            end if;
        end if;
    end process;

    ap_NS_fsm_assign_proc : process (ap_CS_fsm, ap_block_pp0_stage0_subdone, ap_reset_idle_pp0)
    begin
        case ap_CS_fsm is
            when ap_ST_fsm_pp0_stage0 => 
                ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
            when others =>  
                ap_NS_fsm <= "X";
        end case;
    end process;
    ap_CS_fsm_pp0_stage0 <= ap_CS_fsm(0);
        ap_block_pp0_stage0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage0_01001_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_01001 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp143_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp143 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp210_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp210 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp265_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp265 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_subdone_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_subdone <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;

        ap_block_state10_pp0_stage0_iter9 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state10_pp0_stage0_iter9_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state10_pp0_stage0_iter9_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state10_pp0_stage0_iter9_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state1_pp0_stage0_iter0_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call145_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call145 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call211_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call211 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call265_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call265 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;

        ap_block_state2_pp0_stage0_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call265 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_done_assign_proc : process(ap_enable_reg_pp0_iter10, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter10 = ap_const_logic_1))) then 
            ap_done <= ap_const_logic_1;
        else 
            ap_done <= ap_const_logic_0;
        end if; 
    end process;

    ap_enable_pp0 <= (ap_idle_pp0 xor ap_const_logic_1);
    ap_enable_reg_pp0_iter0 <= ap_start;

    ap_idle_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, ap_idle_pp0)
    begin
        if (((ap_start = ap_const_logic_0) and (ap_idle_pp0 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            ap_idle <= ap_const_logic_1;
        else 
            ap_idle <= ap_const_logic_0;
        end if; 
    end process;


    ap_idle_pp0_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_enable_reg_pp0_iter2, ap_enable_reg_pp0_iter3, ap_enable_reg_pp0_iter4, ap_enable_reg_pp0_iter5, ap_enable_reg_pp0_iter6, ap_enable_reg_pp0_iter7, ap_enable_reg_pp0_iter8, ap_enable_reg_pp0_iter9, ap_enable_reg_pp0_iter10)
    begin
        if (((ap_enable_reg_pp0_iter10 = ap_const_logic_0) and (ap_enable_reg_pp0_iter9 = ap_const_logic_0) and (ap_enable_reg_pp0_iter8 = ap_const_logic_0) and (ap_enable_reg_pp0_iter7 = ap_const_logic_0) and (ap_enable_reg_pp0_iter6 = ap_const_logic_0) and (ap_enable_reg_pp0_iter5 = ap_const_logic_0) and (ap_enable_reg_pp0_iter4 = ap_const_logic_0) and (ap_enable_reg_pp0_iter3 = ap_const_logic_0) and (ap_enable_reg_pp0_iter2 = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0))) then 
            ap_idle_pp0 <= ap_const_logic_1;
        else 
            ap_idle_pp0 <= ap_const_logic_0;
        end if; 
    end process;


    ap_idle_pp0_0to9_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_enable_reg_pp0_iter2, ap_enable_reg_pp0_iter3, ap_enable_reg_pp0_iter4, ap_enable_reg_pp0_iter5, ap_enable_reg_pp0_iter6, ap_enable_reg_pp0_iter7, ap_enable_reg_pp0_iter8, ap_enable_reg_pp0_iter9)
    begin
        if (((ap_enable_reg_pp0_iter9 = ap_const_logic_0) and (ap_enable_reg_pp0_iter8 = ap_const_logic_0) and (ap_enable_reg_pp0_iter7 = ap_const_logic_0) and (ap_enable_reg_pp0_iter6 = ap_const_logic_0) and (ap_enable_reg_pp0_iter5 = ap_const_logic_0) and (ap_enable_reg_pp0_iter4 = ap_const_logic_0) and (ap_enable_reg_pp0_iter3 = ap_const_logic_0) and (ap_enable_reg_pp0_iter2 = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0))) then 
            ap_idle_pp0_0to9 <= ap_const_logic_1;
        else 
            ap_idle_pp0_0to9 <= ap_const_logic_0;
        end if; 
    end process;


    ap_ready_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            ap_ready <= ap_const_logic_1;
        else 
            ap_ready <= ap_const_logic_0;
        end if; 
    end process;


    ap_reset_idle_pp0_assign_proc : process(ap_start, ap_idle_pp0_0to9)
    begin
        if (((ap_start = ap_const_logic_0) and (ap_idle_pp0_0to9 = ap_const_logic_1))) then 
            ap_reset_idle_pp0 <= ap_const_logic_1;
        else 
            ap_reset_idle_pp0 <= ap_const_logic_0;
        end if; 
    end process;

    const_size_in_1 <= ap_const_lv16_10;

    const_size_in_1_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter10, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter10 = ap_const_logic_1))) then 
            const_size_in_1_ap_vld <= ap_const_logic_1;
        else 
            const_size_in_1_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    const_size_out_1 <= ap_const_lv16_5;

    const_size_out_1_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter10, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter10 = ap_const_logic_1))) then 
            const_size_out_1_ap_vld <= ap_const_logic_1;
        else 
            const_size_out_1_ap_vld <= ap_const_logic_0;
        end if; 
    end process;


    fc1_input_V_ap_vld_in_sig_assign_proc : process(fc1_input_V_ap_vld, fc1_input_V_ap_vld_preg)
    begin
        if ((fc1_input_V_ap_vld = ap_const_logic_1)) then 
            fc1_input_V_ap_vld_in_sig <= fc1_input_V_ap_vld;
        else 
            fc1_input_V_ap_vld_in_sig <= fc1_input_V_ap_vld_preg;
        end if; 
    end process;


    fc1_input_V_blk_n_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, fc1_input_V_ap_vld, ap_block_pp0_stage0)
    begin
        if (((ap_start = ap_const_logic_1) and (ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0))) then 
            fc1_input_V_blk_n <= fc1_input_V_ap_vld;
        else 
            fc1_input_V_blk_n <= ap_const_logic_1;
        end if; 
    end process;


    fc1_input_V_in_sig_assign_proc : process(fc1_input_V_ap_vld, fc1_input_V, fc1_input_V_preg)
    begin
        if ((fc1_input_V_ap_vld = ap_const_logic_1)) then 
            fc1_input_V_in_sig <= fc1_input_V;
        else 
            fc1_input_V_in_sig <= fc1_input_V_preg;
        end if; 
    end process;


    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp210)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp210) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_191_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp143)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp143) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_123_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp265)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp265))) then 
            grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_ce <= ap_const_logic_1;
        else 
            grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_ce <= ap_const_logic_0;
        end if; 
    end process;

    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_start_reg;
    layer13_out_0_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_0;

    layer13_out_0_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter10, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter10 = ap_const_logic_1))) then 
            layer13_out_0_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_0_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer13_out_1_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_1;

    layer13_out_1_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter10, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter10 = ap_const_logic_1))) then 
            layer13_out_1_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_1_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer13_out_2_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_2;

    layer13_out_2_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter10, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter10 = ap_const_logic_1))) then 
            layer13_out_2_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_2_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer13_out_3_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_3;

    layer13_out_3_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter10, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter10 = ap_const_logic_1))) then 
            layer13_out_3_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_3_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer13_out_4_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_391_ap_return_4;

    layer13_out_4_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter10, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter10 = ap_const_logic_1))) then 
            layer13_out_4_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_4_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

end behav;
2qkdpNPVv4MDNPyYni+NJPTdoz5FroH9mRFIQu/1yL3RyG1qac9899FMoCqW/rGU/FQPLlSkFUkK
v1KMSQ5DOxMbNHMVPqexsbg7fCFyDWn54d5K6U0iNgxyWmobIgA4CJmYjz8l7j3tfRdaZX4pu8x4
+LURbMKMIMw31wzx3TlqSo8pvganzHPUA76vQS6xPXqV0OJAxhcXytg3PSuvsCskKgGwk6TPWWQ5
ftrfqj0FQBpQE0qNaDnLYIxcINQoBRkIMwPlWLbm4NJYKnhgd0ejsr433Mu+zxhJQ11/6uqU6rv3
2f+VnoSZ9wLNjr1CZwYQCIzAshlp11buPzg+Ajhz7U6qcdSqYicH52tc9kDKC8bwz1UoidWMeiS4
YcICfuWXldZTLpbYZhGT+jCeo1Pm96Kp/yv6puedtCWZ1sUmgj+M/mmI6i/3acfmLnQaz9vnec1R
NP62fdTb0QKsbNNxJklF4nyPbcPwhAb4/bcctPTimzkRRHLkN4or/T0TbZYQdC2n+jtxyP1Xqw29
rpVDmrIEN2sriTbt99CEP/MmsUeOA/geICtECwkKZrcNtrmM18OqzqbQ2fiNjKYEZVJ3qBPJCNLk
LmjcPA7rhCWYWTo3Kb8ZqjxWp4yP8/VsCE3X9tR/0r9NuxA+8Lh9TJhhIqqDISiy4iE7qhbjToB+
7WSFL8EZuh8VYdnG9sihKEAqq2zGVHoie3OMmRePjFqxeci1vpPeOw9ttIYHn9JtBojBn5V6j2yw
SYHuV1xp42oxBktxEc1qk0Z+CfiCpfMFT4a5OZLRYIGV4xdGI36O4WrZLKj2ufIS43xWgHiZpg4K
NDXZ757GhbVW1ZY3Bkc29W0YuBu05O8Z89LSDpxRgGu0TJCwMEBm3rhPpZxeHunFD6MuOOUkH28r
c6IJNB2biKiGLZeytJUeFdWAyawGz9PoArLXK4ZA7k0+YifJhjZXPX8HKNlQ+X+NUlMGY5YNag1A
+/csYs25krc3x+dxCEes+rFbyeeu8AFLV4aE/l4eASEh3DusYOCSK2q1A3ihjntuXmGp0f552k1n
7YxlYSxRKBFfeEMARg++fRROsZy6W+VmJjdgX1yg2B35CPhQhF6Dn70NYZI87/rMfv8nDV33+pre
4ik8MQdPS1rwMq7mDJKlmKr78r+NJAbDMGvKChU3cRdkz7HC16jD5I6xljTZ2ayCGX3TZ7RnhDOL
hh3Mg3vGErB16l5XiqqgwJ2Z9DKYq7iyw44Hl5kvMP60sVwzTKXKr4Q9tCPfMxzyFHqvN5mCxycy
gAUdJ8MH3B5Q3z3u3PpcjdAy5gnnH7ntWzTl4hAOoka8KVjY8WSJKmLI0MRf1a/FEzcRI5Ye2FtB
GdyIlz1Zf3ChbvQIkQeoOZ+N3aOUJ/6gefv9SPuoEcZbzQ5KcVAbcacGvQ2CBDZxeJniArCZtUQA
B62vVWulzsyCqrpWyeGQsldD5JsKupENiIvgbtmLeuE8ODFb6tLFYiNAcvBQQ+dymHRMpZhCFC4M
LWZ5k6xGScUKTVgCsphTdC3wmxsu4iQWLbRwe7amXLxhwG3Jpeif95wMMaXhbmBaRINSFLErTZh8
dNyF7iR25jWa2IXGnp0qODnwZbvx7QRsEgdBAoClGeXOGVBjPB1KTT9ft0ATd+QeKgULu9zR9Pf7
IhELgPmwKpRt8QdpLMTW9wK4f7EiKESuLwP8CM/QOjLWUdECncfLsA6hapMGWRfnfinAegfJ2tBm
OqFqnlIpBuql2TxiuvVbDWyevroQxtq7qllPrsKsi6hqPcbScTPjxPWNJAa/k8kCntLzi/zuvUcl
LteKa2f9jqKue1zRsNbonz+CJZGoScsLdtS9kgevq+VTs8kHTCnylG5Hc6ZkcTsYVgOYkUfX5DZ6
1P49T84+ysspZ+sQzLR0WE9K+FDrpIzQcWUzIJuJaqtEAeg+1bcaSg97FF+4b6bUcVAvxtbe6ZHn
qWOPHEB72NnZvIRbhMnJSDi/eMtfZyd45YlUCcsm0BaZ93j1tf4iSeXv6tTJNWlVDSeJ2IlnhYzQ
HBhmxEnObDOyGvjvENoix+xHjVFLDH4fZ5PNGfwR5NoIFjLGPjzW/wpRKBhAjqNIhq7p0UrW8Isb
TgcfS1I9pTzSoP1v/hWKMIAXDDsHKBwSZsNKntZ/yEdG9NubD0/PAEOiEQoQAShKOMo0cpxowB20
YMBUxGNO/lndAbd43K9Jbm9dF1IkeDZ6A8F8t5M6xdUASC7V4/DYPjBGdPBd/AYy6MAiS7QUziEX
Lw7FFGcqr9PpbVlJ5aCRqfUtR8TI9zuv00m5Ntp/Yzy7Icf4hK7YViky9AR61/YaxHEFeZolHJJR
fkZPO2SA4i0X36Yi88ucxH5QVSi88xeYh0njtxyzZxS5rxAHPyI41ReU+Wf3irLjTmh0XBPP2iiR
/mCw8phQP+XpxorJ0j8vRbiolIwPCfFIHBFXab+kz/agLnoyDDYPkf0IxPX6hdrSIfsI53mn1bMI
UzWm5yhPY6EMRVeUF8DSqnKLjIfzImnJbe4Eo+YnPdA1e7eBzVA95/cK9VyUDsEUIm1s0tkbHST+
3W/fWVLoTn4dcTy6QRT7tUBaX+797vcUkANbJSTjEJ358xZvnfV+Zz59UDNa+VJvzKj02MWaYD9J
JG1jIjyLBXV0wbeEmQr2sHBgf3kTt4+dH6Rs35wzJqTVYsz9g8otMJ0xtngDDJlunBf7zl4PkQBy
5qzMSQRbVDq/N5QoaW7z1TTOopI5+cQugOygrI6Tm5uH4ft5EjBSHM8uD3/mjRGIVQAlboMrVYM3
DpJn1cVEiZ5gZ7+9Z/08nnhoe03oilJFsEeRAcPYxmUgzsRBLyHhHj+C8EvV9lVzh0jPCBm2PS90
6Dj+7uR1GqMMzQoqcBkKf72DbREVGAa01nra9KfmcXQEzTbYIgFKHoMBHjLaKgofHR8ykGupxOqB
b43ZtJpAHJ39VRBq42bhaqe5NOaRwQvGV8DROmVQh7pPKpBdfjppQhygqNqV/KSG6rqKzDNwiPGc
QCV68IgHYY/621yroMwy0zN9di7zQ8IdxKg0iRdrZqV1GdXvow+mLDRrsh2z9LrmHVwpQk56JgGW
+wSAgQy6zxS1ZwzWLO5Cve2stbD3to4ADVStlOtKGttAf6GN3dlUbso5TsshW4EAL+CXt8Pmo+Ax
YwOk+4+HznTjInG5dDpss+xpgxtbcTnCCaWlky6dbweajlo3qeu4215SNbwuDgXBl81CT6J3uZyO
aJg91h5BwXf2TAr5reOLLLKyxRScjWVmEPuki1YTLM9PnbJa80Oh1pHDWsdIqydNubiREEnOScpP
BE7GKbd3QLaF4+XPGaRKM39JIVB97CH3ueiggzN5Mg2rprv4VtoYKzjibQ+LHJ4uPvYjAcJYpShd
pHJxal3GZl0XRDD/rCttsrypXUPzLLhdtmtzRyu9D0E5HsuSCG2mWDDwIs+SVZtYC1BKGwc63c54
ucrfGwfWSDRb6j7o+OKLQjYbO5+tzUQShPWGvcLgR9Tj7zxa/JUHknzchk7EvWHMxG8lovk7Nplh
SJuJMydNm+tLschriHwDKFMr2QdNS44e/ijZE8BqrC5dtjcUTSNYuQC44K5HHs/hSlt+KBLriztQ
IqGGi5v6s/Zburukbmz8s2K7DdIFmJykOg1PDz5k+Ajk8K1N59ySN/UNWc28A553fUmk5VzlgbpX
YE1DBryKJHEddUdLdk99hFRVr6UFD/PjOxg5GLoqnjz3PGVVu3Zn5rEdpfuOkGBxm2228NI1eTYU
dwxmeZKeYSYzYZTo3FM5mDLpt4ggD+qgvbWjePYE5m+SwZZC2Nmd2eUpP7EOtDhKwsl/bwmzGZ3i
iDmCcAVkwtTAIn790pGA0N4f/t10BH8FMKuN/SBZnmfpJSpcmu2iQ2Uz3u1Pyb7/eyrfbjN8Pq7Q
jbBCdf5dsShXS+WFs0Gc+KQWHQSKF2KbwXQTkfECXTrj/qsUaNNwi4cEVzUIQRipuztd8YKNjyC+
+8b58AnAn64oVfp6rNrx6M1fF2CvDtFqrVAPJ/ARRY/kiJp9ikJLNPgpsvihTMfSvBCnW8p8COoK
16PVjuYFJDvACqGhekMDOZI+pqvpkdeQgV3oZ2TfwURy163LoBz1f8iGfYRGk3uQlXptcbOHZTzy
+xnTbcc1RDAR57cOcRsKBA00t0BoTFonLkhehpgo5eAgUzp0/mH5DJ/RKwZ6qYXvfATbbXUHDhf+
oBVid4MsmvvEEWuCS9WODK2Hcn0EE2f4EcCqYpjczJGxeEWTmkyBZDof0v2vmNfUgyU3N7qtHEmN
CgwPus1QnquXfnRaSX0ZojyMQ4i3oIwqXRBe8U0HtjTGjcNxYqpBTnlDQRen53iQVwRq9jOOIKmD
N6EtFXzu/U1l2B0vWcugfjh5foV1bAUpVT0xNdkxOsPI7HpnsxWdXfBKUUGZAWTNbPjVv3QjIZym
aLBTirsGD0OMFv1m4ljF7py+C0wuYyDk0cNBgLuzO/ci75ViZdfR/cUV0810ZEyL/9cKh/A633WA
hSo3UJcHsKbduwW+1IaKgHfY+Te0C3JHJ3zhB57wVbOqG1QMbpEU8f5x+yqXmHvOvnExJTgTpueA
IuapbonUNp6hyMd4af9yBlnMfzSZMDCNPV7nUH4dzXB5ctOFQrwU6g2Z+MNECYdQTphuWrQFHG+R
tKzdQyz9Y6N6LAUbCEp4NOCZu0w9OuNSeI34RGLOr3+IqY3y6+hzztXGvfy/YSa08E4CbPwtsgON
ADi2rh2Oyp4TLlx+Eg+DYK6K5E67Z7YK3ZKctIWTRQ19Ju9/msaUkRYvnV/0mHhTsatGJoF7/FFo
gPBJBq+JymCp7UJiE9O5IGXjZp1sopw1w/LSF6xfkPANB4yOGcT1pvMP0dYez939um0II9SvZtaf
PcCdxQnBB9F/41jrUPwmF0zovPhSnPrP78UjbVjoxOM2iwPAX3o4YSN5RJ+oVWiQ8BrM3YaDa/Fz
00xzOjzyzQ5kQCudUb2eTqfIrjMdXmEmt5Q6uR8MIj4cUhB8fUMKMZCFqrNsuJ+lHtUJrdFS3PwA
gdEv9jb3335ESs3hTFwPg4/142ZfQPVMlU6sQNi+gJSKLwqcL3J/KXYHLRjadbk/famcQxwVlswI
JFvyaRRG3ATk/ueQdJ/zEZErIFXqtQgRxzYFlJInc+bLaD6rJf2yXUtbA88eGNEHFfutc0H77Lv3
jJ+IdpFAWBV+9Py7miEizf6xNL6AqKNwES+Qrl2h3uaLqvgZgd5Ffr67QnUDMFSi3mLhc4pfIA4l
8Ly7gwHRa70muEXCK1AdTqaiWheDYO7D8KGcZ5NPhSEuhqOA0z2mHhEyss5X5OMMFk11CQG0PCSC
ifXhvd46zE7+lFUSXXb2f4H0Zuv2UC07Kb/j4VMHSkQ6AxwbVR3HUlq1AQSVkag4sfLCsGwILObp
mcAbFh4jOSNvZaPCh42GwftHBAd5vP7KGXqQ2snxKu85MsSEpMNdHybazdN+07CUsffov+pmdadQ
ZxtEuW63aXQSqhMiW9whuGsZ9itBDCOg9W98yUeb/T7+F0ILbnUS1pxT7JJzN1pP2ZN9dzhVuOG4
vCsSvFVxebAIcfuyZxIvII4sLqh99okfcwvc1XENVKFcO18N4hdO2K8Oel42uHu1YYSIvUIb4uqN
GXPIOL1XkYTB308ETMEhpCPo2nZuEqya4uofLnM2F1zy/GSViYFz0QEHyhtVYrEdEjwsxiGVHz+F
XVTzXUxged8n3Dc8NjDV+w15kD4fTsyiM4tnwz4NK9n91hf7YcptdgqgY3Pbr8nS3qUK9e5R9Yh9
mcGEJeZMUHRducuQoYSAQyZcFEX2WZ9vaBxW/FqNWOUrvtvjxOg4l1YzsZCHSwn61xfeyOnvIUcw
NJrqzS8QIoyo4rmDxqySyYnsfPtGCq4fcP7GtMgPzo7aLhaZunPmNfwhyt5Z3IkpTbeZTYzwzNP8
b7jhtJ8fcR/3p0Q7OpKpE1vqgIP+LJj/kh7wCPb4wulDDvonqAo27ZSuP1aDoR5yblzfwg3GMOpp
1yxIwekyjeorcIXW0am2s5ZsRJ7Yyd2cLqYd3CV3FyVIhEQ/+tYecG7r6iplx21L48lkg5phcDrb
IAGDDRDFxBPQPu/MhpsiCRQjz+tQ8kt/X5M2a4z98wj6wCl++zaXxoSwAEgSyVe7zPUjoyxn20X2
rG2emGLJS1zWRO1ewGXaTX5BKAsgGCFRYnqrIU99+9Ep3hHq5A/BquifnMf9pstVokN9gy9cBpD7
wr9Cb8JGPv5KN0AHtXVJR2Asbb/wDzLxRJWIh52A5fH36cQDgtOQTJaNfBcn7Ckh+79RMFcPjGYt
N/IdcZ/J4w1jNJmuHsqq+k5FcI3+/qWhfQnP4ndjWna7qKFyISYYmJkT7VgKFbzDHAwwaRwKuFpv
CxMorL5RCcDckgI4nYwT35o+dLqI9Lfo9hPyQmkidykCMfXVDpgVIxok69Pap2LcErBBfwl3N+sx
WCIuk+wol7DGhWlesfwAvz/B28xGvhab/54HPU850bkFZsFfVZ1+PzvFOXQRtM/UmUOwI2V/OEYY
4Jg3V9cv64HD0GKdwUut5vADST7XAXJNqvVrqFwVzLt+9bMRy5HfPLhUCQOHF/ln5aol4LWVGe09
k4kzT/tWK6deBEfh4zYZ4UMaeQZNuLzjwneqKTyhU68lrZ0yht8Erk/PQeqV8o+8jDPwFae4fT/b
JDKonpRw/vYCyWnOEhaZiqWIkR2tdgXgNE5dWAHB3hQUImVFJ4ajgCDCGqGpuVarIrU2SVvXZggE
aUUWrpiRMwvyDsAw/6OnenQvO/gf71aFVkwFQY+sq7IsViBcFunHdYqURnO2STztQgAP49dUnTzM
y3i7wyMmdS7yrrKT7xyTnDb0oCHyVG7yHYdZtLkEbHoBQvnfvB0lXuZ2AlrGPWk/0j4skETwFTWo
RNrQzzW3Kwz4FmZtrDYWOgMTlcZ3DLGgguBP0NYp3gWUn3KR3HtGEqXOZwZEXRSO2nR04dt0LGX9
9K6krM10N8LcQ8O/fbzvZqdTfP/xUYU3NFAtOV/r7dcyPZjPloPYhaUYS31aDD9NU6v3ZBpwtiC/
yEX2Z0MylCa/SEByhpr1SeCHwC7n5kH/14yo28zHgd5+QDIUm+NMLSeICmJJIFBBw/ByT8omtlub
7iKHCbGHbl0OZR6gs575wLj/q4rqcprWa+t2MCLZYA0Ep4p+vRwmN8VJCFInLQwH112GuYe9RYn1
VbG/91jsdcmNhnAiGRB+76lwBJ2TUCivrQLLw3GCv7WytybBmxve222ismPChl72U+tCQeiHh4M3
eloBa/kmIip5jTf2SEGaSwNB8qtRwk5GIR4R7ICsJwZ+/VoZZp4XGmtxGIPUD7Fy+kLkZ24y7tLe
pd4hYsKaSYmw4tHW2yW5CxnSiOZnS0qoE5E6VvlIT08Qmz4jA4pEwswwzwWZ/cUOxL/quf8gEXeT
6/N953HiafU5Kj9ZSyuCfiS1a8Mm2ttgWYiO3IwhJRedlSQwbUMp/3BfGpovSKYeFRPHUMD1scoL
HKuNMrYQnye0lMZ/FltA9bARob2GcqNThvA9MqXIwSICZDkx6agx00TF/Fv6oVz2KaZco9KYk9Ff
HRrZLtDY9tHpigaS9KoIOUjCqOHCcFAO01hKki+xpG22Ipn1ka6CZVeuM5E0nJv/9tP1opPjDYEa
gAqrtuCT8yAMcRCNDYTu6AtPvsaxMu4O8A3u+TxxEArvv+WlCYl+EjCGT71O8x7MwMu3VFSG7rC4
BHqsWSEDDopcalMgmz8VP/albSoYY76W5Y/vzGelOJlhODoG64hgPM7fLF8JmzWv48jOIXn7WjUc
v6LeeizRD1OSIbDaDbKZHqg4lMUx0p/dGXiT+QMY+RwByRmxLUeUiCbhBCJAqiTvUDjc5uNkoHhM
aq/W+XfdiEPch/0ikPTGKouYTppxex2ZFWA+/VdjjAulh3Svm7a+S2F2yfcjNzNHomTjrRUEK6x2
je0TKFSGXK2xoB3BAkRtUWw6dA7YtjRg2SFrzuXOXT4V945ZPzSnJOmjdNdh446Tl/BH0hUD+Esc
+Ezc2/xKt3oD8aau7w6B71zjpA63oojKbBl0/PN5CcRjGGqlS9z5r4GzkSbNaND3UQ0c9SzXNzO+
6qgSrs/j5//E/VxArg8QTE6wgl2sDbYiaUSFslA1ppwGl8Rn6b4SzhnmklR+zFyi/AC6AF8u350o
CBc8ftDa5ZNVXrnApX7RJCtMYNK0cczEWLTjRBRLfO+uZ38tTZ6VfQbBs2GG+sdPo55+yxwbn9aV
GVnB1Ogyb/1SYVITEh7r6aeMF1rrmkYQRDHfoCFdYmxompCLMY8CaVgC/pxqbxCixUk9GKp5qwN5
KeAMTcXNtv+Of3lD/CoYMYcxwxS7+AFUe9Bia2tFvOsYGxuubpEoXGz9JGK+R0+G5SIhihBe2ehq
Zc9qrRZQ3nW2O3p2V/26Y2XApoSkvoc+/qscjDxAxGIIrTmwHZxZ184EK/gUUW+D9D/F6FbNmUfP
l7ETnrl/6o9EmZIEvc+D66dJ+bOry098Ptz9Lg6AxSiD8idpV7dTkyfZAdeeVKzjZuTzxoBcSM57
Z+gu8mLg/P2APojNeMszy8fV2p1FkLbj8ee1D9Bd39Vt5XBKcqUqDxxr9XOPfET5ml3UUjkQbgfa
u37av32KVZdvoX2pR8wpUYGSTOH5/4SuV3JrwvNhJCp5HeG4yRYF3+hmPsVBQToy6jGu886gb8FO
h2a4kxQ7UP6Jhvfh3aleyXjaPtRWfxiwRx/i0TmABI5sW72WFVsJsRvbn15Od6q2lwpYBF1PoarE
nv/pQ1T+n3H5PATyP+YEtX0DrnctcZt00sRuDihTnmjVGDzGJUhsjdcxSFPvkVeqf5BWIeQp0V6r
KYDeWsbyKlUJRw96vmR+5uefm2uGJU5D5lL6DHxRs05z9FCdYuYVwwLlIMaUxbUiP+Mwpp0pJMg9
YEkhR9ZOvlizlaqGrVgg/E60GHogilg+dd23k44lEsmOtEr8FxHwQGXTIyTQLjodGMx32GyPnDUe
csmiBJuCMptKzQaukckt7fKZQBYGtZc0irVN6iNEqEVPFGQsDQNBrUlTX4VOgt5Q7/XEo4fY/hK3
GPO4fbmOop/Ss+aibvkWZFREvWKINQBu5jv2WA/69cM8K+/fHUx6unkVz7eldb4kPr2eh11NBr0I
aF2Q+PdhZfSdRCjFsNq4J9iK/wsdgpxCAbSD0vTrvGgtNPGzWsy2jPnsNkTEBnk/FyBC9o/o7p3A
p4eMwlyhNwf1hPdr8IISFOY7ckgadUWb+FpPNyg7FgC8VrWupv1faMG1fIlW01X8J38ofqoS8bZ+
R1JCHAwatX6ElcG5jNr+MvdpwsKDKIx6dJu+mqcJdU9fpsTlATHxMd8xzzUO7fJ10pogUzZd6Uem
Yro7Y1K0JInpW3OKJHxlakCiDbUnrPKPrJI1GTLq6P6x1qekA4Nz0pFyjL3+in5CKrvWyNZyYXik
x9jjG1Hy00lt7fjf3VNTC72SydUraxzTXKMcZ4UhzYDyTRINHnnLtQEdIV7BpDbJgPrcAgE2Uxh8
TTkMt3iDspKys6BrcZ8yZkYp/Lo+aB7k6jLpL+6y3uMMai8Xr5jqwD5zY0Ei5+zjMK5z8d+XVtqp
xDa1MOZ/CKqAFf8SgYOKLcH8BenKpLflQYGLpwnJgt0pJjVm1IPfUDVaIjlPXZKVJckuIf1o0sUh
v8SAh+93898swVZpqq0kPmB7+EFCsd/rixcEBrd4IqT4ZX5Aaqd00JmLxkUCqB3cm4pTXcPreRb9
LdyGZ7hx57PodfiJP1+9AbDxTLn0hKTMIjfk/lMjdryyFx3Dyo8FT7odIugmpMVotAtuvuZQYu+Y
0ZMUec4FJLut+cvaI3TvkWTgcUzYvudKk4t3K+POuxdNr34B9+51sGbUNzggDjd66YefbEeKPCXc
tfD+Fl0R6JzxLFHgT5Xm882CB8D4u9BSuuvd6xFNMOUbZZhPWzSIpzYuvz7YUJJamHnfYmDVissg
t3wv8RRR7MmLsK0QoZZEXOl3CUUYFPgyfUZHaaKG5veauJzoldkXvqzRtQRYvfOvaLHTXPTHGTLe
qy1/1o5da+hsTdPUMIJyLCKnQ15fkN9xicFX9Yft82QqjRVWG/Wc7x/ubze5DYHB6t4Qb6Fxfhuq
urLP4spMujM2dmI8zvKC+UiPvFEdOr3l3mPoRcCScFEtRFqvBUwPhtiD+bxvyVcc/tNkWi1sWvv/
rF0g60KtIq9ke18/LY6fTp3j9OayC4Tchxjmvtafd0uA0HkqTlp0LsMPK0Pyf1Icb0ea/7HProft
fC8rq/mBAcful7zhhf+PfHwXD3AxQDc5dFzAJElSYvqAuxVBc9ZKoRxhdda+lbO8bpfsbuHIEzIu
x4uHgXUllcDfV0z6Lq59v7m5dFMX2zFP7zcCQZoliEDwyxymM+GIyyPyTr3zvuXH8vp5w0GPmWAo
215S01uPfpv++PJSaGP7UjqFCbUtGTzS1gmWk3f/+kplq66hizhwidn3WijHiA0Rn1Mwgro7BmfQ
E3QfyU83+JCeYQIDcmmPZRimOzzJ2gXGBT0LKzt/rswhyRKKARqlDcWlnxkVQFDkR2aokB86+vPH
mNF2QQU2ZAPr1i6Q4GURIhxd+KHLSE40oWyAtmkkfMkKd4VuGguUGbku9ekkpPXKBng6DCXRREm2
GdsAVujoAVbW6TOwnV43qqNTah+yNBqCh/XARo5WKZY/Pa1ZG8hhakfqvpMgvRIOtUglRbbIdQJc
Q7kZO7PI0yL226PIs7MlqBkoXuVnU4uK6BnjJjTCdXuJr2aX1ULTXoGIHw1jNNDotFuNTQIZS4Ai
HVXbuyCOpfoCROZGEe///rPZWJvIwJp7qriPc92aQbXGGY8zKfVWyPhgDUueMGYGVcvT1/CGDQ5K
bPbjU5k34zP0s0a6jIQII7DeiZUPQHPDVHqUKGHHze+FcjBucb0nG5oErUHkVWUexgHd+gnR9KNR
p+fOnooG+vG1LPLTOXz10TEtW5Y3pStyytIvsPNl/KgijMLdmwEATB7tVy90pIchagqPSNuCOvX8
5ubdm8sBzUmK2ouLjaUoBD0Vtnujp43CWIfVHuf49IaFz5YkDC1odFHQyEIoz+MIQz9VyTRLVchD
y7L+0cvI17IvrJyo5QG1ucBOsDyLEZO50VeKkeYFi2rtPIDc1FyWoMR4bTUk6HtayBPglKWhB5Ci
nP73qcOYzRlrtBj1kzGbRxYbN4Ja0VwGwwQ78mzF3galIWBI8pHhzc3iXZlUT5v36hLPelLx06vB
BmPQ6Vth0qeIbY59mGhqRFn1y4cnLrRz22qtTEd98AvpQzmpm1rghLUWmKFRm6o4beevlqV53Hcv
RkLbkg70YSX7gSnz0oALnamddPceXMffXuhLU93RTd27yxaNJG4j1u6umcXS6DyspLiQDjRCE5oD
v+CF7tfWHXFI7b6/IT4xIpYWfU1TK0zHPDaCTROHYr5kCDXnISt3oFzbMCDkRd020Z+UIfZsoB8D
nRosyU9sgvDiRfN8ec3LFbdG6xL4ehBDWx+LRhj3Fk+am5MmNPBzq3nEI9yhwFf0kdVzy+7Onckc
q7uMEfh+Gz+qfnSWQCUsx/vRAVhO3CSqvxI5R0Nsn5AbZm58IrH6ODmE2jGgbf0sZPbFgOv3UnWs
mOZxVPSK5AE5+syNKQ2OOatrJ1F1tyzC3WhSdXNxCjUjqa01RH+Kh8MN2iakERlBs4nC3e0ScKUw
QZn4LvzfQTpKbucV6V5AZiD4ygmeWQy0Ex8dWaY1wELbYItGTaE2GbWWU9f3OYPbeBAqJfj3gcdM
fr4JoqGWM9VnWPL4kwntGYlcvWKXzQJHp5nGUL/vi0dThgr0+BujyWM4l4+nn+5/JPqre80TIvB+
zu6TjPlTWlH7OzeeEHLOf1G9xQ0gDFy8Y8dJ1J4fpKXoAj0G/3Hl7f9adMhJs/Wpjx7VjkVIKVP3
G08LcrwhMwX9m83b6Kqw/Oldpq7mkIJy6ZGjWENCXnoamkHbP8E8LrxZedWSrDQxElvSAEHIHM6O
x9+iFULchiLRObmGn7/2k11rjz4n0DN6eY+VoFBZ3pL+j7JYiyzw5K86PPVcjzmg42SrqHWXjVJF
Kg/VNXPbU6dHd+dxdjyy0yUz19il0B151vYZVyDGEbHUN/DClWMlo3Hg/VE7la5H19VJ+4Sj22Xr
P9tIwt4eh9BA/Ey7Bsdz+A7ewW/mg7RX4lMZ/YMx1ou8VLn4IK1v5lQ/M/4be9ZN50dfFGUBkNL3
k5+fopkQT+C6uXyJIr/tHUkmD4VT0eHUfUR90+IWyQD45AE2TznkIqh5zx4XZk7gNFOtGTU6QbDn
fZaLjXXwc2kzc6GVDqvk1PSeMjwUlsQ3lOAKEA002OJKIkZ7w7VSIcXgIK70+UCQAxWAC/3JEVPH
0m6qIxJmBq4XmHQTbEloA1/20Q3cBK/U1gMHSVefWZp0kQjKK8PK+QTSZOm59jxtIYSqjex0834p
iCRAIXiQynUuX57I3GN8u+6CUjvthtlebUxIYI9kYicd5NIe1h1Xkf9fp01cEFHazo1CsNjGNY0L
7pRsMBZ6yEMRaNiELihSL/XqkNXBN5mMSpRPQrEDKyuZLIMK6ZAs++/yZ536NrOf561PcrHQ8iGS
F4zdKu617eAxWz2cPd414ivPajRfHuQVO7CSFWTDh80bDG2rj5CjAZJdWTng2+S9slitnYZ+ub8B
c8hcTAPk5UWPAqUBSVRPFkHa0mDS10fjvwiGY8m2meOBxVZsHfzGB4UU8gdBSAK3x1X5tQ7zFIaj
aVN0SR9QtPSkoyjI9rpZ5rj2cGJuHublJgmxxnasQ+LjDkjuC1HFexGZ/DIn+/7O2eAF0vgZJvRq
dH0Imtlt4WPS6xqClZqhrRHLVbhtxCMpHwBkw6ubYfEXtz9MEM8E6UURsL/oclVocQxhV4NjMiMp
4XXbCcl1BPxVIdct+Ujvx6MYfKu1DyjyifledyAJUrVO6lsUtdfeZX1ezcYWyHBKEdPkMEDYczwA
yfKzIkp+3VsXwtqr1YM07z8diA4fPfIyv7nyjFfIC3oGasjT+EUJgJwB2lygwkOJ9MAZeparlEss
FCFeC2opWgSLC60V/NDdO/EOm+BtTXLR29MBDWbFSu7QUCJA8pLpjo59TyrSIUSGUtBv9MCd28kU
7f9Dk0WU7Bv8ZmJwM8nibG6gOVZNpIWeK1F/bqdVaeVLpVzfcf6+tLGpk01nq2H3KmtwgWTX+WJ3
0G8+PnkKjH4BILGKh9FSu3Q6VGTvUQlzVhr/82oQzOuLclZT6bzgilwQYtDHgRxMrr64mjtdWkJf
9cnlA9RbUaVTBdjC/6K6Kq0IebQzvimBnhZtosgxbEB5W5/k0lZGpJgYanfxg+zrYXeQZsTMVIHW
uNwf9qusxv7peOtFcFl/nA6xgo5HEOzK47EukrDrQsPKTt8TPPTq/PQx9rVJ05reAMjl34bD/A9h
Z6aDsUZob0VRLRpw04Dmpr0H8FSrdFQRLt5ghHW4rFhuJvAJMvgFyh4hxmHHnYq44SiP60s7++r6
XPyOKlRmWOzDdlii7JX6gFMPp1Y8PpixYo46DBXAcu08x2ytVr5PKTO6fkWjjMUPe6w89PU+lifs
MlO8x6HpRlLYjkV/BLwvsOTbXks8I47Py46yljMM8qDheisqVIx4QaJHqV9PJ9x39MSftosmjdEE
a6yKaBwFsSnH+603rK70AqAwg0YmXIIFxnnYYKxrVqrNSosbQYmm9L+O35Ax2M+mbLgqVCfcc3+B
0ormpsNJAuI+1whtBaEPJl8h/jxqT5Brk/AtuG8mpd+unZ09A6MjQ2I7yv69OBFwBl3cV0IQyuko
fgl88dOqoCRjBXiIX6T0u12/v0kT3gWscX3sZWS1pPaQnPweg6foP1W2f8Wqnh//rHiCd9GgXE2H
h3e4Q0YM0AX7cyk9Mtc4fw37Cm5CpGXi3jcZ/aU0tZK1moxjxO4TXLrG2DgenZHSKlfPjYEb9+mo
Ocf2IWSFZEPC8Lo0JJ2F4J2/d3rYRwTAiQpfCL29fcWKVnD4BK5SrkWHqFWlchpAeu9TkhMXQQbt
fHUnOgKhC/n/hohfyCv0fWvdptfNS/VyXp7404SuEAXp6qYXYHMpjixvom3C2r45cnimw/+h+n47
EdpFykhU47B8Tefknj41wbwENiZ+q3XL3m6siM3iy01pkZYMKL4+yzPEGjmbFPfDEh/QuVlQTEUE
jvy7RF2o1fZZn3mvy2GCpcFPPmYLzEdHHrgHPBJbiuM+q5Vi5hL6sp3jBb3cW3/Cw5ibRXHykadZ
e2JyUMlbTfaS3l+219tee9Imt6Fa8bgnbOmGrInN9Pzm1pdVtU7FnGjAOFIaaklrunjR3Tcn+/0/
iRnP19vfuoaEe+3nPEjRheRBCroj4AHrT/5fWbNgYtOEjN3xRBafdkq/OqZfdqxYm5oCjJw44RUZ
ETfZtVaCD7xuXGOaIpN8DbKnhDobbeHE+1m5wL6VY1auR5Y54r5kMNIcRLVYNH9gDyk0ccMyqbP7
AZIw3UU9Kd/ps/giTwMz+bujXVNI5uY2bvcwv64p7d+ALIVdUTqxMZV76Nn0ZgGfaWNGWOYIrSaT
HqqT8a4CJKWRx8IQSPPaqHpJ4xrEcllo+LJIiqk503+Wr8kv8pDZQSif30wVaidbhDHi2gG9FR46
r/LbjAaA7KOF/ONNv3O1mITaglvew59tR+mlaEE0emTbctwQJtLmtFiPNzb2u+L+yinOEbayq3Aw
UI+IxiMYId64HdM+hzHuJFZiPHG422CSxGMLegDZTrwZ4YERQaLlVmYa5XyvpYTofhy3NRFU1C4x
lGd/HkSqVM1RgsJsbqIxR1OeKxdbq2ntS3gjEX5gzrQvqJNzSWzkcRwa3RjvSVe/MeLv0/0TLbEy
gz0/TMikLLu/v5B/2lg68EBmje047SI0SugnAVQcmJGIqvRR07RKW0Jw4Vtd/DKJ7RIKQcbLa5zf
m7Ay1GwrVNtAid/6mBdWUjhRrQF8gpD/pQbZfScjRj02S8+T151yWZeG6suGWLmPkDy9Q1sUWJHb
dho9ZGPUHPwdDxcbkzep5EO0rXlUJ5/yOHIep7bSoJ9qIeTv3JKZyPKOMS7cIyhaV6uy+e0/M0/N
aigQH0t9HABIDfyWD2wrU1P+9PICh1Q+1MGqeiEpxhtT/f+JDlVQZW/NG6+g5Cx5HGtPlaJ0ogEs
OENr7XHwgAeG2f7sZOrlHNpmWox3dzXWVMfsHeFY7oVKVhMTeWAAphwgbAJ/Ozw+xWr/3yXNMvPO
5EJm9vo5HFUw0aFeftIbFNrMhqqrXsqvyKkxGSpeGRa1WsWMYynphmjZ6AQ61yF2uW91OeOjwzzu
3+shxuL9c7QK5c+eP0tT4hMrAVP0/nn3pRRWiR1wlibXlIL+blDPtACPIITGjGfu5fkB/N9hwE90
AYrzODXzSsS8V5s4UtczDJdAossyT6ruvYT2AZrdDZ8COhf27E8q+yftBOU3crcndJnxCihoUYS7
X049SRvAgfwk/JHZJCbOlJJDsr7ggPJEKMPJFNiYExBoocTN6Jl1/AhLSIhdaeiQT4PZHFtvSvzM
N01FcbtknarTsOk1Qbiio8GTvsbvkOgc6AvZcZ63C3+Tfv2aPxqhSBDH123beflidPFhQd50CQu9
F0cR+NHWpmr8jIn8EAfs8y2ToHhJnPBINisHC2NHAyY6BOxxQaJIflAgIGrxZNQAiw5pfHP6onVj
uYPpEqSiqvTD4r248RFhWXGrEzyiRZNGchKk7UEKmXoKnalgc2V0klPe1opVqudmBS97LsazcNkF
xZJtfHzpIBJKYpluSdds4wui71tk5hTanm0h4ENSlCwIFxOndSfjEZulqotKb6vIBPHtCaTL6Mwg
VUjdUIICBDS93XMfNXS/9MCb+59sBSzAQkOHcoLxO+aeHvEivN9/0EqDmkjUypQ8/ap0kTJn80N4
wZ9O3ypoSIdbezlks1lt4w2+qCs2lpht9BbV0tyJJPIbS/OTdM9qF50cSAZ1DlEPmoRNZeePt6Jy
GEJ+43Dsz8P/KbUJW59Q43wR0KOpPtMN1SaDXlNoxaJWiSTLRrTAHcH2N6bfy0+Bq19TJsj3px+K
tPQnPFVoS0nosI99MmjtbVUAaP1rNGePJBuxn5pvPNKF5Ks5RknMbnG+Hn/bkweDbmeeYK8DWILN
QuPV4D4hd621wiGSKO4Fk5CdNcV6eGT00CmEDXsVmlcG/0xj8KuhW7w8s7vkTi7Lv2CrBbz2Rf3T
VpJjA6hqKNm/bsOFbNqs2vCGinCqr3Ps1Q/g+6jDXLnDx9fENRYZZkNcgX0gLzWteo23BmUI4U9j
5vRlp8lLNhzpfQkVdH+uqVcZ30YOCx2MLRJZ1N1weYnmomNO4iMXeHqvvcFRxYwb5FZjmQ+0Jacd
YQMHLTauoPIXoRYk0nRl+aiLIAX0SlGhQ2lTG9KqWMc0IkrAZg/WonRRtHcThWWsS4Oi9eLUGJ/T
c2/Bi07UQJuYkIJeVenWorII/tCJV2lmB29YpfVDxbYe21tsEmIRFptll5bYL03BSlfps9iVaEFZ
BJMsR7/4g2sxUWC+FX5nt+L+1TiPmbmN6M+gQ73ZEh77c+rGXRfP0OX9VM69qOPrelGCUHJ6hYO8
RjjPhpYZTE9WvA3ZN+JZONEkQBLVN8oCmCSM8AoQxqZfnvZ1zg2v4UryMBPCNdg8u/JuqJWOEpCV
12EE297SzuSDVuyXTHgKgeEWAM0iRNkigGLuU8YXZh4lIYBH0Bua+b1fi7aaTCTNjD0OLQsblQOf
aWu7M3gLqPt+Sw8VhPk2DUXQmtN0Y/WOXKG7k4rOK1OYqR9PerY1PfnoL5Tl/9mUG8McGnigEIOq
94WrYxJ8twjZHWSYBXZUt9GTcgZZrIZQtXpY7ScrtgXeTH8TjUucsp/9wvm0zFB0UiDTpxmGLrZM
c+gCY1dvlKhLwic20cVXYFVASyg6SXyDAUSpghMKvew0AcVTMJaenhAQdqUeDpZq9wQo4mnyLacV
Vq4qcIOmHhBhfIaRH+NdYYNPtrWBPdm9wx6QT14bVaLy8dkYzkSf8pt7qMOfoC+cvIxURsuVchgN
/To7gUA1vHsh+oaChFRl3211Uhupu/+kaiWgE0kA+p39VW2iHuv/ONl7inx9JqFhoHZ35H+f+g/c
UKRA59/r8RdMsyKI3xu8cU1jmqJLgMT5PpWfFlHRLEji8Gd33nLL3fFuLBKJONSpUJnkMDAjnUne
ys7moWLcUH0UhVOu11hUAKXP+CNmEhdkxYu4NJIppaxkILj7S3bux25augPxYBCwPzb8n5+3xir7
rH3sYrp52nHAFzROcnszyfal2T4qzZ9wS8u4huxA+TaCcZdz4CwmpMw/7R0VZb+JedJUrKSM7BRL
ybEL1y8wc0aZ7efoSd4nLW80MJDRxztcHdLv94QNwuoLKogk5sDxOLiomD26uoTZ1Sh6AHxn3k13
B0U7Ub1YR7Do0Wx4VPnUdpqKbEhkG9nhIURRowHCLEEbDf7OUlvIbV1O8yP6CXZE5bReRPX4d4Fk
8CHSAdCKlbFbkDSpAS+xLkij0UjUPELECRyxn5CGQqhoEEE2zDGwet5sJnk52eVRDSkA0VN6+PcI
wThqCTFC5WXOimjdnGlF1UNVxoE1xH91PlneyffKdyRrBBkltdib8DYWxgAzA4pjsZLjgyf3X9Gg
/lWhkftv14s/5PnwZtn9GqT2eIZeUx20eAjQoXJWEmmy2EX7uFmh3D0j/OakyT+j2XmVGEQzX6OP
1ADzubWmj34ik+VSKku8+5X85Wdf9/dNKuBynJd3IAxli/5uLfWTFQ+bfVqM+fUcFrdQfPSgc7tU
5wjvL+xK5lW9GEw3oeHnlQ2loHs47RmY2InSQ+z4NYrGCGhoMBgmNjv3u0HYlBKdb6EAG7mJaZuI
/VZTWa7PT/LuRBGdNR6eJVQf0kHBvfCEL0snrgeNSKskeqCtK8q67r+mPujvMcSu9JnKNCOpbI6k
AS5Jc2QTYYZ/092j7L2U+SVoQgK0ch/N+IU53p0cg7j9eEUHMDAJHobZ2u0EDVd0gu1DwS7x/EAG
aqInis+7zgXwbgEvjX5uuy0nwug8AjdyeqeTWMcFHVutObMNVvYIcfltoS8KotmPgTs9+X5Mkypw
Lh+h/QzQHWthJ9myRiW7ysGMAd/sGo7V2V9/THBUOQ1zxjR2GyH2SfjbK9gBKOTx7q5t0so9yWn0
LUSGjOAaIV8VRdwFHVWR5BLUE5YJOymSbJZ2dQ0TMjVKJ2fmohy1f0E/n3ExZkTw4wobHQW/7iPa
uxe9oAOiPyIePGNau5T3QpkCGu0nx8NwiWNb0Dwn1h08yFsgwQOf77kp2e74vCrkW3kIh/Pisu+k
q+G/wJC9pw9HnFRCWwXnlfjl8G4gfgeWOWjxCpX3DgoOf5/1KHG0B6VyZ2S89jX3ARALovXJccPt
2K02GMXXPuFxC8MRELM1Dpr5oba5Fvm99kF5wTOWvuqX2OC7tmEWdANZNfOuSTb0utiK2e56QiaM
KTGL3tChdf09SFb+c84PKBfu/4GraPKBtwSSPdMxqgm/6Iyw1/p8/mRFrVfHHUsOo1KtNHl7pNFf
tOQbYxr6o8Bo3BA0ne5cT2Hhu/mtD6IK7wL+2nK+DR+wV6Wa86qd0QYOeSRLCoJXTbOxqtdb8mbw
ErovyNpAWfY8Ha1YilCRE4yn+//rdAeomxcomYQwJ18vW7ATReyOUw0SPdAS3eFdufyesHlntEw2
bqyxTBiosOOfxCQzs+B5q5BvClSazIn6K6UdQdIjXdqayiR4nND7/krZmspjBSJJrMrNkav7SSfl
d99xPFm4RSkQC8FPg8ujnRsH1JCx06wthU6AcDgi8if0qHIdgeyIOlN14oJ6NcLL6NKJw4G1CSbl
vYJD/kZAaAmaXAOIL9fS5wwYGHnsrcgnIIpqhFaLJm3u3pUPxxxetIZBw7UkBPAJTqYH9ejj50AO
UvnFaVZubnQAQfq8y3ebx6FEpHv7+ni+LuNyPdZoNs2HHEqsatadAL23JqdiG8rR96Cg0/qtXTqS
PYvZ23fqOeL8ohIRF5YETYLIEfyOWgETbwcyJG9yf/5bKALoxKymBV+fKn19l8TwPf93FUsQVQgh
tSubcbCFTLDFxMLoyRssNv03fYUinmfAtyd9C5VAYmJJIXry4I7pqRgrKNiV6MdOQ2LJAquN3jfM
5drA24N/8RpH9TEsUtlGgozjAazxbuYkOl22yy7AhOXp2DuKXyPSUVmgbFq8Jik9vf3GU0x17k9n
5HxvEtHGWtTOpozrYxDOF9P6IQ6efPkJ2jLWhUm3smjhJ9uMwoZkGfTrXP/tEhiZErO5MOcRKtQK
YupMovgBF8PaNklTcUJ0MVfVh/+fAIeHycE3TbaVoxm9TfpOfOqkrDC2L1jWZNF/xEp7xuVVsfzc
BSvHtdVNexbq2buBrbix9f9duyFmc0x0ZOjBrsqiOZDFOVf0XIuCBbV5Hp7hokqzY3i7kqB2JxpD
me5aRvNU6lwIN9lNjBdEzojSwiT4WV8O3QahKfOQD4fLuXnWNMYPUagthOekwTm/MoYSZaXotWJO
+cQBeNazve48cigXzZVeVSRCjfC31tnUd62uueh9QJTkU5dBpN4P8IbK2ijV0kbCpgzDaueK0gMF
I9TxuN3g+o0GUkhH6xiMYRT3ylUrBCff/oJHod5i5isVyJmyA5k5cc/Nf9Zai0kiy/4HPRRKed1w
qsKDRNwmYU7wjtf3rFEPCvTbi14IQSYFPsvY7HO4SS82Mn4zJxABDBJ9fcBcYYWZHg1wjku4wbi+
LIEVsWQt/PZvyzvqcztgGRv8GL2e0y38WrPWhZHfGuMRjiBqJTHvyOB3f2VthVAcUpnbbQmgDHru
aIrU0ZwFQGHU9r7ya0/ieeW7+8LF2En/ZZt3K6as/K99SVRJEPcV/1KpXlcwLBzLtVgFmFtpxFhg
Mw7wH0Y//qoRRjpi6FpK98Gkv8POWssgFCf/NUGqo5QcDUhdpQQcj4WbRAIugxVIbVP27XKRyq0m
Ms/DYlcc/sRQ/MOcyz4n4h7zRU7a2OF7F5imqfOQPG4AYnfTB8ug/DUEqe/eV06gealw9o/qzNGm
i7tIud4D6G98tzfFGNvPGGxAE0VuVkIn2m3MqwyrHljVU8guz4NP3Yu2Qxyb7W2ITjayJ2ag4yMM
VBXdW3CRdG+hyhb+XEM31o1OBdBuMnMR2Svcm04dUbH0fxOWCZM7ySAxnYJyTI+ssP+8RT/3y6Gw
GG3WcOsdTVaItrz7kAijCeLkYsDXqnDowRbS2sddv37RIUnqwuBqIv5IL4z7rxoRL7dNKdmAUqe9
DVsTh/uzpqwmiSuWDJs1CFC/lLdxYAA6tYpzEma1ArDoM0N3UA9Cii5yOqDxx1eTfO/Ec6cZmfnB
Oflg+u691G3ZkpKuq8lMRvghBNVBcFPlXZavzP/QG/DdBXTM4aLQVaxHXtqToWZR6cECYzB/9ZBc
shHyj8ZjlI8WLHELee3Kq8TwiVSoogUtE6rkt+ccVe9NkNwFyJpUGbBYQ2fmUxWHY/Rbj1sRZj77
X7dolnU1737XPG1YHJlxSGCij5vx8678T4qAm0GLK+HMowmJ4X70jjE6fRfLBYgAm/wNpzHVREk2
iGkD38Lt0MkqLJpTza4rinAgKrWwkWYGL+r8y6C3u4HomXeTQtAHwhOBsFAPcZ6/8SB1ZSoOa2xs
LcX7OLfHe/OuOuVHHEUZwhdgAxfwoaG8ShsvbFA4iMyup2fVBnOkPIgVaJB6Da7OdSgltqhOHq1M
DClzTxF8XALb9CKwV+PsAAHTK4JLSMoX8jWDqm1XVg2puS7Sh7WTN9CPvc547R9RhFPIz1Cj42oq
7rlJvZs22p5j59+9Xnvs2e/qrNGMXqLZxORgeYqvMcov7W4Jy8YlZJY8izQHv8sjTKWYCBiu8PWV
RWu3VArFSGpwfTVU4S6SHo0dFW1S5lgXbJmPlipBzjGddWG8Xp/sG2zgjf4eDhOnQNiHpVOdLNrd
7qQHyb0jhsWDTi4Uk3yHtmCuTzqRHSkwF/XwclGxQeUSoy4GIv955wq0oSLrcuaeDJcoFWgixI73
8gWm5L0ssxl4Pes++GUmakvMMVnVCYaZ5WZzyhzcA2v8pWLSoQo4/tdpG0wmNWCMy6b0e8cPjtzp
A9WCsmDpasNeaGG031y0yLZdKNm1FViUjPaadknz/B5qW8OzRpVsAJInhpJcMIec99RNyy8Q3Iq8
LZGV7xuAUYmcY/VIuCn5PAI8WKI8U+BvLaYm8pc4SpYNZE7yw22+CsQPtoCrKXpUSEUX/ZcZ6+3P
jJy1vE8LwXxr4dI9gH+66991LM2ibc3s7z6ip9I+hM23X29uZZIcJaaLXKtGo2RdmMEuRRnsjrvW
8eL4g4g7kk4mJIXiINnsXn9sTPP9uRAQhx1MbvDGGnSPaMh7RNs1ndas3pF147bkhveLcYAMdkX8
wx6ctnbqFZt/BxBZp1dgZPeIXImIwb6lWYB3LITsnkO+QbDCfdVeAEbSOo2nv2fjkwGAZbHx+VxS
IRhTD4N3Id0JEtJZEteiE4WNb/t3w6bX0H5L5L01LdSfxaEBK2mQjoUBnvOo/LsfzhUHdh2Gaz0d
cGxwDsoKr6MhOeYjPWab0BHtyaj3HAlvjnaW8RcpqFAUwN4EcGoh8j5RlongSRRZT9KfBcYYblBI
7R96iRCmZTKjB+d2P8bii3XhKiA+NEj8OYrKUQUIoDWQ8k36/NKa+TGf4NDpxNRlOPpUutHCRTzl
Yh30z6LoMfiMuquInvnrJ4SdRFaz/Bwb13OVbQLpG0N+ePQKibGuX1W34uOLsKjVoHh3oapoMh8u
BTYfo00hiYprMUdDphQXFKtZDgFcRa74qCq2O0nVb/ndOlSuKem7dnVe9riDhBtLuX0J01vaj5Tr
mcNpjZ1H3GRVCvyX9KvtkysAi5pUBkoZvPV10LEurJOOV+K8ikKkdVrArb9GwBcoEavvI+YEno/z
a9ql86J3tonUphsda3oHfr7xJWdRO+AlKQjCf39E7QZ/RFXQKtANEgkxuD/vBsmCi4TAfPrpOWyC
Cd5hCtpzqmr9kX+CrVpJ/iWxaEmJfYrLOhZp3wKm/anuz2f2BQrGS2DRWPyi/ymM3bmJkfXZr827
Ipmf08/bIihiYe6RFZE5p8UC+JSNz/EPOEU8UsUyk83toRsXP7rqbTtAsRAwijk8B99VUWisRSyq
+O7mZ1EoX/cRvZExMFolgqESgckPETRrSSTn85L/VubL/hie3fC6EBwY9QJfV13K9xlkIspdygqI
rJcR2KH03/739+qmhwCC8m6KHm8EkmElfRqqCcB3k6Vlz6Y7Pb4AWvES4AnNolN/UqLLhUnPgouS
KK/QFngSVGDvTGvjA3HsZF77dxIADalVahQcA/lWhl/sXkM2IxVFO/c/fFsykO+QNtu/eaSYLfR/
PFdl8K8CSFpyrc3weOiy+9ONpOXqdL+y4v3KMhQIIMrSuDcyLffDLzAePl7hJ8Neo6AHLAObadGp
Ht7f58pf+fCLyTBIqpQHWiz2/g7MPQ9q6HuDWb4LXLccxQQCRrKijMizFj7CiwLAh1SD0A6OgT+g
yRHeX97Otptpm1J32h7HyovOGQ9/0HKSOOJ2jMK/vLb/fHGDbbIaASQMd9WKooHNyIwjmSFfLD8Y
KEqvbgv7fTFWVT1lbZW5XLwuj1IhvHok2ZoJyWj5Fs9zuK/w+5E3m3wHFIwg64SImGPQRIrb9/YO
mcFGWclgt1T7Px9PhcQqccurXxrjiWXufBXjZ9jkr3k0jgzgmeEJltBSGw16ADF76TEpGXkF5C08
IJHQcZJQ9v0p9IWpRXAq+fY1BxSekSn0FVBnrS5Jf3obDiGpCVG+kJfXcsnuv9nJ2Ir3BruNwXTG
1DDPvNNbTB3yFPr6ru4QPNfPVtGjn6iv3OsztlJjc+1EQnh31Gufqk5MuqV/+Ofycu1OhGX9aOA1
pZn1AfzRqHNLdkgxmOMoCv3+xRivRXxUZJVsBHVzkL33OjxyC36lfRLuaykpT1GCqJ3q0ijcYqLj
+e7y4QMN7AGNk+EUsks1hs4dDsKndpgOC9C0KoTc28Wiv0NdYqdBhUBAWAoF5SpRBvz2ZrbZw7Nd
fQTotBRxydC3u8mGmbW8UZq71cPchfhDL70+nwFcHZg5j414PFo9lodKsBRdsd8M+bRr4tvlcYL8
C80gdESXOA6Sppnkj8xmyWHLep8j6ThI28Auv7nwY1m4KdgVdsu8TaU+k0PeMYdput+EQDA9eqwE
W1HvWwANSTcNGc+ny97yXADV4Gq0msqk4esH9ONVpzNB0jjQGPHTXwIFvEJAK+XRLDKZ0Yj4sUaF
Zmiiq9wnypwOYQ5fJ2rqQ09apBXoS4BO59wdHv2uD7QvzSTI60Tn4IhxWnJ859cbztNCuTh45qk4
AJC1cmnNf3/XyS93cUfQipHjtNRR+SnO/gSgqHlzAy/gLreHWmuxV1/NNSj4iUouB4M2hnh9xDCC
mL/yQBJpHFbWebTPKcCYcrh72kYzIwpu8ToBm+AdxfAreWoQCdNnGpehEM2L40gSraHUISJg9djN
IC0rutknpb6tMW4ckRd4ySD7TVlClVYtpYcoYvkWWhyxY2hryLIsw20TP5quM1cjD8gcIKcPJo1j
vefiw7HlE7SeAySz4RLgz+d6cbfZquqlF9qs0J7VmqmcTfHoXfB+2KmvTVR+k2hVIx9klOyo1ETT
XrRao4AnmBLupTyif4zL4kWa2X4KymtvFxySznTUpb0Qvr08g6ehlc5+sMulSEXR4KzJNUjpEwvs
sWNqE1x67oupHlJCeUXm4bpQSM4pWldloI5+MBV8TjHlusgeWSgF7dvLgDU31px52KbECtsKmaFk
b+8tH+rw1Fx6ID+cqkvqIuqsejjQ5jNGC4nmWvNZk2kgEbrZkkDGO5Rs7dsZNepd0Bcr00phyond
vEQi04nDVnqDc1DWAmv66rNwkA6BHCCviRwbnAPw9H1x3BaOPIE0ErPlZL+RAN7hdikoYelqDIC/
au2RLTRnuW0LhwIiwKigexmMPWnXhlQyqx33VOkhmeOtDtHi1BLRP8eq48QK8ZDTytWdYxU04Qzs
Hy/nRqddP15Fw/fIOx7V3G2vJrrNLE74dA4rum8gsMuykye3QYLPGdwUq/AxpT5z9jD4NTZFiQn5
OmY2Kn477UqWv7esX1DfZeTInq24igJqhP8w9YKCZwdvUdQw4TJskgCHMkYKWukhQ5YbXcPCVXhA
DY7pTYC8ANT0PUsqKtWNkFylXrHrz9MfR/jUAEN/Py5RTjY2M69XeisifgDWPAe4V5Yr8yxaWFcf
zTzY6ctfNTyBIhTR2MSqGx+bhfTRSbkEnT36qoprsb13YlcwVUHMz8ZR6KRHvwW0pIppMEFxWmpf
8ZceM0/96p+qjkzu6dSsxQSnPpvoy6p+yKanEPOqzmr+TEdeW4c4iRFqSakmDK/6mtv+WMlCc2Q1
wyLwqWUsjv7HMT9KordqrRkm2TaYIzeAQGhvJUbMJak5k6ofMGeRk3+4O6WogCw8kzLOdrwQD8mv
SiZhBdNjSUUT+FyJ60HbJ35gBl+Wt6YayP8L78MiDILmjL0m5A2FSUpCWf2dIVi+GRdKJJo9uk07
bfTb1tZwXd7ejsy+8IQEjjQJb+M3b76N6d1JNKmIFlV/K90adcKCqxfiZiBnGPDwFowMPmRWpzcP
0Lz6EUktIvl4mAQB01n1QUSl1Sh7C4ds4hIBerSlndT1cOs3FOHuojWkGlG4pOtf9KoVFsRXN7GN
NUqeJPdQdxlFSfsY/Kn0Ln+duBtSLHEJYhLj8bMUH7uN42p5RjIqsUhhbIyvmF1txT8s9sJH/9f4
5l7mMGj6tO2Jfnfkr3clCGnvfS+qc7jVL6pvLpYJSI6WHR4MlCP9qioBiE4u7jQsT1WH4rxwg19Z
xhm6xvzcU+AfMjb5i/mCRHveJEDxTzU7rkcYHdryu/Jl6JG68oCUDg+oVU9l6PdUmfkmsv61bIK+
d5wBhiOJJ/sdSydd3QXjDFb85UnffHLIVT0dy/+3uxNzzcGMKaWlsKE8cKkkz17E/VlWjd+VuR0e
uM8jMogkMZmf+gn+6eAFskiWuorAOt5P22nbglBe8obuhC+L2mhbJNpcOrqfp1evnXDzta6LiACM
FXYQk0lhAtyH3/7uT7714TfMaS7oSr8tgDdaa7b3TzPaSJsw+xPSdDfj24hHbVTiUfA+Y48SZXGF
wSJvU+0tAGWhLnzwOgZfV2OvE1Fq4BUfq1VTJb/00rW24SlDo3OiOY3IbZE7fFX7gXGjmWUDzgCh
14cPyv6cw5zoegT1d5VSjaWKNPH21gfN0WMTaQSmBpSZZwpzQxzyuLzY1QnhiK42Y3Ybd6lRuiTp
FuqCgqGxLiMmHGGWXAj12RGEBTgrelQC8eZRWaJvIZPIgdVf7MhwZ0/ReO3lDD3FxnFq0q+5JA8S
Yc+Kri3rNA8BcrrLyjvW+cJV1GZymtIlbp6VZsHiTuvZHTlmTVKNUmG7pBuEM4e/brkNmk4BSAuE
Nh6wSfoUoI9skM3YCjF9tlkMM7x6UfqI9d22bx6Fu6KcGkmfzACDNusR2dK41aP6VRuJOM/y082P
4gsC/gH1n9A0LrW1dfWq+/jXVWbSoxpfor1s+z7sXBstRRHmKdmqHAEkcqsN9sdFKV3zpaXjJ54e
ADDY5h2tK0XtWAuEfjHSKSx2mTqLAtEW6Qn9V6BDYUKMECrFbsvDgoax2KushtqqB+ZMkCNjWHjP
65QTgbu9QLtad8hXcfPWlg2d6yn2a34p56qnQA61gmMEcD3wcT5xUNEZp21cDEC7VZq5JVgTQP4Z
WM9WKPfjqF1oaGnse4Hglp3221J9f/h8sKOQ25+UnkHpnzkshUICFcLwhz9z+t/FOkhRQax2S3Xm
61m9Ww5syMAbVk+NG5QR3Ty5TStqqsLitmQ72EvgY22Chlqz9GjLf94BWHHmeoGl49L5oYGGE9Ug
c48y+OIY/Jrt5r/rG6BmxEJ56g4y43VlumOyLB5QZCjAbAj9M0io1TTr6MEDaC0z4H9yNCifyoA9
5FOEGBQjDDAQqp7TjCj3kXdwvJKPfz+PGHWrJ0qPKHBgAm57jH3iXMZVZ7ILuucbwXP7+gPWs8vl
CIucm0b3VFATzppPqwyCnFKgO42d20HmsuF2VOzI2fTP/fHzLVZrrQL0ESZSwlOJRiNpix/CxGyM
SoltmPAPXkpoi+SlYqlvIMpu+qR0JVy1l3jdOQIHYcMqor66QlkRDsAL9BzfSHSNNxZftbIQ36YV
3XvYViSDJn+SwoH+uwJVYXp/kevVsunKETbPGZtP01peRK+pUlnbZWVetpsej4jUuiBSdfzgrKUf
6KDWB/vqktpNqc3kLaBl7X2XtiqEyBllqOdH8Vscf7HiyERl40pLxgFRxwZntvJiciVxSdBwUOfa
denqm+fzOq48rzeAPp4MODkIbswybO4f3xfBL9zg4tq9kEO0SA+ael8jPuGg4FEhdSr5/N7HWn4c
4lWTadVJj3yI9lj7elfoadaFgQ75hoysFztzBQEnwyLURlRmx0R3RBzaL+wfaVOtBJKg1ssNLKzv
PduY/BYDrSZDfUJZ9EyipW9FZN2IXS06OdfInE2p50RXx9tKBT08dNx5fxknGEHTw3sWPSJy6r/q
8wO+5qT+1SovmsExJeoG2elJN7zrsX9gAy9xKMoANaV7o+9JBuAu8BB6fIh+ktmRk8yR1UTsQR0J
G4492VlCBETHldEi/jKKWT4luZNcvNsiDxPXRe5qMeujrTIK2DIt2hz6Ws/m+rRYMLCwhBYCeUSr
YAHD+zsotvFGIUTjBSvxRIyiFsCxZFHXkNwwRQ1ovFtj1/n/k7HtMG+ijU/Y//g6CfB+ChFkDcsY
Mb/txbPN41cvGhyXQsVrONOBU8UPCCPfNqASz8qv2dKCy2SlgPaAtRq3O3EZfJw3Lmb7dZUIoxS6
MoqjFWmVe3Z5vt7aowBPECVrh3Fg0/rC5Xrrn2La6dx57KNYK97VKFPAobB+dRoFIQZmZBG7guXt
prNX8TQRpphCqvQ/vYQMQkjaq1RbcSq0tsSGuSP1Y2viZavvVuyzgmN5QvpVVOOyyav7w6jwZsRp
GGkltBBUJ3ycGwMBkn+eUNYLrvKlV2egLc7/PaUIk2IxtWjCd7qXKGk9XUyPwND+PTxtMvzwf6mj
39CGBH79prxluqj6pj8K32w6l/pCXEP26cQP/obanXXhzGFrRFZSnljrf74FcWcChVQ3xJ3XafPH
K2bDlVbnl15HneWw51LsvibsHq34XXnM3cFUixCT9vXyLyKbjH0msnQwCFXYIAZrGudd6Z6OK9aN
u+WP61oEOc3UBl89r19O6nbd8ik8rszqRXXuXxYop7YtiE5oAJk5Th6kZhqcapUCbwXC/pPnOKdR
QZbPEyZNeA4/XWNcdRbwkUUGlVpVNsi8Dw9yow7WS1CLuDiYfSL1o8EveorM/uSJRoMbYX8V/wia
D/A2ridIGDuXA5lLbtlBnQSb9oyAOWnMwIV47oFlLSDVC7feiAslJWYL4jcElIhx2/Ydvm8XXSsb
9GwvIiBPmroi1EQj2yC1w2NVZeescT5rB2AmLsIbQboK9L9wp/doh2aU8INaiIWqDmOG7g6oEMUq
D3hLOISetA84F+0t4DYu4U9tUgvx6FGwKnTz8PVB8K13DTTPtrXuGnfShmrIRaxXo9v4ThR4XGiF
4/qBHIA6PNdkvacKs3aR9JzS/HSDvmUQ/Vrp2IO92vZ0GmRvS87wvzw+Ap4IXzdlmVoH42BUqqTL
IS/8Xl/8re9mEsYEN+oJeHvBLx/l+Ggp5545GZ5Mn/187U5F1ouWwll6olpjdAfyqjFF1kiGO/2t
HbRvWrqoikBpJj+tzBupcMG6mG2TXybSQv4S6TMC6jRNhkjLjAXvXL9CDgXaxMpcFxr+4OZnIj8/
6/AdoKHMqFPb9OjpKYVvPwmtNi4e90VJH7RV7pU/k6p7ZkhqvF1GTbjDRqiHDbTTgpl+9vjRaEjw
yn/Eom9aeRMKylw/jRi9EWaHeFtO520TI8lhMuCkJ5t6gUteyqw1clNXyyW8FDbkPwQFtix/moAQ
DVrILyWtcREjU+1dbfiw3x6vbw4GJVSRz+9WN1AaVImVSN4YFC4xscYzvXreOhpxI87K9oDGr1II
tVeMirm2lRX3H6Sg0EZrPCgjU/CwPxfL+R7E/j92P0PESQQeHi85dp8fytSYY0AgPy72oYCr/wCP
BpTtFxoGtCScToUYiJ4id3bYwHTlxZU+denEP3jGbfmWL9S72n6ehk01+BqAmpdWoDbgIXo7EG8J
zApdGIbWFr9qtCQ0uya5a/StP/RQHBwgZP//vMFbSQ+NJW6dAOVbs7l5PUeZ5VgSGWTsouMDbTlM
bQQDaYkQS4vEXXieiR3ezCHPJhjKp5EkxAu+WF95gY0BS6Pyj+3IGYVRC4XjKp819NiheCig9AJp
7LBlaEV+/rrtvznrCMTxU1W26FfYWKKqu4nusu6lDExjmi2sjjowUK0Zzs9aSTQlTarPAoRALEMB
YqSO+Vva73HRp469uy5Bs21VGs0gEJ8igTHO6eD0gszE1tYgt3PIU06C7cvdW3niml4/zomXGCLX
BDLfgbpyHOdn//mIuPxlQOlkmXQF36Zx8yaoIBGlahKJHe0u6MlTes97Xx8ieK1FZXFXtnXghKcI
0pc1gBnI8lNS2Zh7v5WFjdjAju6/IrY9ALi2a0m/TnMOWMUXe+Nf10j96fWAQpgF8FfmMC1gWy4D
TsIY2tJzGCDVJWOaIts+c1g/ZwaoCJ+oGQB3ySjbtj+EIMPN8kNtfysyegl2bhh+k8jZp9sE3bJl
1Z0w+zhkBhWzM2w7xfIffhVwJkjGUewwK88tXh7mh/gr8rIzdqCU4fS0G99yf2YWqapNpeDIcogV
nTNe8l8goR97hJKgDvvGbkWwNJ4RgyizwBeGSG+DJ4wtNtT5THReM/q7xxVvnXOp5CiaOEUWWaSE
O3tzGdU/YFyyI1frQCi+RIlgpbfSDbOfcrTmzokEamYm2fReeY8/g/ALxyzd8ALYyTn4JgbYu3Q/
kcjqZkDf0uU8HV9v/OGEjdxIeKj9Drp0nvIB/u3yCn+8Oe2OQleVRWN2mgXbeuy5vIIDLTOM5fkz
sA2+rvk1+EbnKG1Ge2p4x/BXPBKTnikR/5iBv8EOBUhyu3m4BlUVd65PQcqbDUB/7Of7RvQEBACt
YCYylk9JlswHfYxJV4TcoR4YJKKYHeBCp8xVeJYFzEKQ/l6tYIk+Aa9aCPj8fQEuVt4ebV4dlnco
M/0ZPLg422fvQJ+yj1m9SIdcmgd4vDDnXW6+mN5BQ+VG7PYMrT732dXLH33KDUEbjrl7lqhJEAoO
uZZrXKAPFHMi4FEazWqSl5gtIA0sm2ksm2aIE9XGP2J+M4EzpFI8KbOkybjXmijI0CtxOJ6r4ED3
n56LTzS8IUsl3twWy4uymf/H8h16X+KaX9z8b/QVy7q2O9ngsuVGaqB5TnKNWMxDWDBg/I1ylW/B
MDVmnvawgyzaylaWUHFwRZ3ggJOv/ro0486oYGPR4BqEjSBuQk8C5LO4a88OnnciXMYwm95IRiZy
IT4z/RpvIY0FSL00orjg/wxNSydiyZrkNzsZ0S2m53KZ4YGcy2vaXU9dRHtCvXu0DVihQz/20Mg3
FSitIuY5klFg56O3mY8BSZo7NTlHiZgkYWV8QSk8vysjO/8IGhNc3SEAl7J65o2V4RK1JSwbHl/a
Br1Hp2W+8SPQ5X3oIbM7HlK6C0q+8OTYKE/KhcLjaTxYslv/eeqFmxRHKGS2iPMCfup3/PgriokF
90eSDStTzdaB6k6eUmu/QsI/38cLFyk6iSFZPiJ3qfySI5EWbEjCXELFAfDMjEGCktiQYkLdqSXq
h3CDnsA3ChVsxyWS0A5gELmOIGA0luzeD1G3srY1y3enn1TrNqEt/fCglmpFwOQr+Yd+y7GHQjVd
HLdvg/qtvNnDG1pQab/Jeg9Aub3FvTF93pK4n1k2z93sVLxBpIL9Rq2n4C4PFK4tVP5boEfT6NYH
BdgBz5+RifZ4KUWho/ZZ7l4uHeL95gg0hr7imfHBEFi67MS+eX7HDtTw0zRiYDsJrW+iS1JgPvIh
H87mu2mns8LQ0qXQUykYwUtAR01X5UtnHhAEfqBXtZNQDkkmJ5pmcTKjhqte8rWjSu6W/xD+gPet
gyfdLL4Y8gr3EllZsW6kZQpFr+YrzNJ1Yjan4fwyjhQhjtleSoPCpS5RePtRlLDB/gNxf+Mwjy2k
qcd0ev/WkklO9t8tQu0g/Zrtqr3txZeH1C2/5PbsZxUjrhIKjcWgARpLhIsGEf89hcptP2H5qbvg
LyJG7gwCL9QCgAt/1uiY/IhrKQjFceob5K3rFlpJf6rE/Zw3l0JiEoHg9735vXKKWL95gkDKAD7N
0OupM5hp2w12rqRyYtVIpwWstotNMwLiy6f0IF5eRr0jH96YsomlIe4N4ScN/8qAqIQnniqhwSBI
xIjh5YmQxF8P0Z1fM6Z8TQvB7eLmYAvcdm07Pp1WZcy9eJDeCunqTtzpqrNZvmtA1609HaXL2LAM
w0j7bkugief6S0PvRoEJfj+vYSmlNPS44NiuYmGE7dsURp34+ansmTJ9SZYycVKADjOSsAfiOA7X
tIFvrOOlRawPV+9aIIKlmNkRTLY+ljYQHKm5vVfwCgxCYPjUwtIDYYukT/sK9Nkqc3LkHnOK9YtJ
t0SmnctiUimRjY1o/N6iGlTIR394Mqeipm1zB1xJIln0B9FQiD3rLdUyT5+KwKJYnID/Ra2WUlWC
PrbIyPGXsTgaYIaZXfpxZrYLc1hXrd6qedeI7mDYSPygDtQ5rFD5Lesdu3eD55welcWdZk+j6tH4
rEUg5GurU0bTZwO7mbUz8lJI3aAhiESkolT4AOGol4xbWdm/02MsH7uXxO+1zvnP5d9HbWiGjAcA
lDBkO6n80Bsj5grUyk4skFdyqckV3PgquAkjjjv4aJRBNdQFcENGuMxsFsmsfDnSAZFTBRMyGC+N
UFMnUPmOU6QF/M2Sk8fE7VWrp9jAMQJaJrEmdLvOcDy41htAdiH8aqk83Sxn8N1EYLg6nJGs/yND
JkDfBFw8c+RRHy7GW24312c55JRhtiy7mDMxaD1UcD9NmfvQO1j3oF8zvC+CVvsm61i1J5jhW5hj
TJtpSih3Ma0xUOa6Pu7wh+zPwzG/TXgOsqhMlcNlrGbXJYdlxXfOBWnozyopseuSwlOWzlTvUiKP
69m/gWXdBMa9k05fVyjiStxF9h6hXrmnh3cCDoYN8NEzuz3LPAXnUWtCFbBeX1ZMV4+ey5b2buSy
mlcCKnhJ3Vn+bNwx+YTeTAqXPdfwedw1u7oR+6nsOKI1JRHgxGO2ikyqmPq0QHPlEviffKpmztTA
NNFkdmbDMh0a/CtGTN5Zvit0VKlYXzNm5KKFba9bIdXEHfh+um5+wtPhdTinRSnX7w4GLh6AiA0A
gbbB2atXJZQnQFgL6/YuTbds1TQ6hfpQsN9+Hc+7XNP2rs4Ou8ze4FJNSTu6pVNdeCVwbKeVYSFH
uRyQDcGoBKOXQ9OGrDHTeMvLyXbF0GxNlRxQ0OWQbI/Jgj3er2myoG8/uBpW2+JnKHTJWSvlzZa6
ywCLLXx1rrPSeShhLBxNoQpZxbncVKQBHJV1Tk2q8/2QQzef4sTeLl8R/VZRBKYRi+6GoN1SHiO/
mNy3nLaGkcgB0nOxbPfFDWaDiEVXtVQTZLW3c37JuneKn/HRF90cJVuSrmNS9UgObnl0O7STys98
beVY3jqU6MG0RjalNQQs7Jw0U61FzRZr5oIgg5kYDCHr+cijQWB2J/8cDrs69rmpKtbmZCxzHXiW
qeQqkv8uVgaXzRX9im+Qy0j7lXmObv+wTyvdl5Co5Gdg8hFh3ZzVqD5W2ASDeBYv0WEThBuPwQWF
S3VjS32Y9FRF1Dc37JmT0XjlFQL+oogU2g+xMRuBsLA9w9QSPOIAs5xCEqeOdMfl1dgT5QA4N2gc
yLe3jDohlTvPaiUtjttij7bzPa86PV9q/SoYCUJ+DY13DAlaPhokWFhUry/vvblM9ysxd8lYbcQM
IwMm33CAKAAaUYM/qgsAcc0ZLVTvCUCKmSF9mE+RToFlpD0oU76RR69Y0mchw0ajoQGXy1bYvzb6
shX9iuUwMT4uTmoJpn4VUNt9b9rXiDKsvpj/AY3L2wW6hwx7TTLw0VCPTCLnftRiiH9MNXmZR4bm
Wrx9YvMnCGsQ1YSLAPXvKg0cTg8ohhRy9HvQa0qqwD9B7DCfiUtKf88ZjydYluQhbPm9xcH/S6kv
M6zlOEPLufJxsEWaNm1VYTa/5NZQ47UGKV28KrQdtitwBHWZaHxpuYpObT9ppeSUFywPjLt95648
hPum9ktrxt6w/Uy6qHc0rW+Ol6YQqLIN/uZsyPw6m43uhWAmVDgzpfanku4LrQHVqJXHG+I18y52
pn9q6dUnI/n2A7dJPdxnfNZLWKRMKf8m2rQloadWmjsRBmx+va9EQ0eNOVgR3F/WBaxF/Uxyc/0N
ukyQBFVVL/prpo/Vk4axDH9c+4jBxVMl+bjLEP0RRRNZqBV7asnvupa7cxoHx2E/Ncfar1CpiXyx
7yFExs53BO+NYHwhdWGRm3GsT5Z8qN40+ahY8xSvoMhFVLCFgyXwwV+RPWphAWSzE4ic1lTf03rJ
Tmn2d+1tk2/NgMQRIfLrV1rsUxnmtTZT/NdAG67FlJUhn/ahv9mwvCnY0RDiuo73j5oZXXP2uxzv
rdF5lDYeFv/PNhbUEbRrsRlkZs87yLeBZN5zyLN3lIK6yrEcuXju6HAuxxNEKKbXuBJlzXPid1Eo
3Ks3u7Cj2AdIQBNlFU6A1mh6vjeL7lmPKiHs8oApQCNKvttvU8Jm/8tgnxwOvwIqz3CYXFwrzCvq
wBeLBESik4pUb/NUSDoQiySQakbI1kXPLNMqK4ChLNXrxHZKdmbRvsuk2BINdoCnHIuRZtDFmgKj
kbVYh+hAv+sFD7TO2YjnE4Pz8EUyMjc1bmwyMxnfontXcGo6BowFnp7EhUzcSN25BCXGTAx8Ynns
A77kwrcAiHl6NQ71S7CY9vM6wWFX2DKXHIJ7tGGmaoFOPU0r8UL60L7OjBB6DnDtKxF4tCdqqr6b
