xH3yJZjFS8oIvpTVoj+ROuWsqZhassgyd0CWqxTV8fDoSHbut43VIpFRajLDVzn2R+32xCCIEVoV
sakTH/CgsSH0cb4IG7DmmmoVPqo9juPG63wjf4fQuE91FuqbQhudgNkNI8eJJRjQHhHjFcRYPZ+t
kcfaQbATaKAsiA2kEAk/SCRNxuH6XVN85ZqJyRkrurfOB1QxBgHVxu/vPh1d65yO4t91tFLwABh+
0EXiyN0wk4yK2GYt00aw3TGajo1l8UETtGpSGuD760bS4Op9TYR6vFPlNs8lA7LNicxrRtfNxePX
3CznRKOzyC+m1+eyUb4C3+H8AF5YrHoqaADBJEB5LdAhSPbdvkJ+fXaI8U2yRMXZR9hIJA1xtCG1
qolAhe23P10SWvt6mG39dxo0s5TGruf4S7/0wckkT7Ur2hDh45VcsypCKDCQ8CXD72AKvE9i4sSJ
vGBUgnPJ8yCg6rd/1jXpYWsEMdET5PCZveVaSd6Oxz6Z3HREzIs8iS3fh/DonM7u1j3BjLjbHtva
R5rK+rT0YCi947CdqokED+rooZgoUx3K4dx+pO6xUZvrVB77PRoP3mxnW9YSwAPX9eBw40Qm6M87
PLHfbQW/BPtPtoLLiTS57AtMKXqA6WOpBxVOxnDO8QQ2tyBCS+mvNcmY8ZY1h3AvSF9eg+hm+pvt
fpRzyo0u8kwiNU8hF1KDkULe22vOSfZ7TMW+kaycf5AJGcTTfwRDqXVQPbXcLSzq7E7yS+fdsdke
6Qd9vcWc2RQe88hnGil+Jrbz9rsEbk0cckDPwV9AJP9v2B+aWKil7dMkUUjH/X4hnbVJIWb01pQm
5OG8MXoCN4mhv1fBdyf+se5fmaOSBPuyJSD8MXGqVfZYy6YWmxnEbgqtHbs91eo2d3hJYx59e8N2
ymB4j4O6oBmjXFJBjkVmHMKBLhXAKcXvog5MME5slPywc6kgMZ7VsAjsCJETUN6aecpqNjwVIyM0
ty1RM6SaqPJAPEEORs9e+OWHgQA1za+H2BoDZD8gNOVuNMhK+WZmKboLUlahvyLJC7JNXgsxw+Qq
lvBScOfiKki7q9XXu8C4wlWsGYXTtLB9fhqyDp8eByzKCmsnuDOUZRYXACtUtkva2qtPq4kTeOYj
LBR4tyO0YUqKNkU3TTsMsw6MLEQTGVfVN04cFUK28JFpoiwfcyDxt6k2EHfGsr5BUZCEfzoJQj7l
RHeuZX+yEyGG+NJrtuZVG71SO9EDCrv1ckBolcwkfqO/G+jH1fFoEzK4p1J+7P5JT8LqsKhIk6Vw
ZqksdmNwar1iPayCylaprf1+2qyudIsH/7GcVB5ayxf215Bf9+Jjd+pKW8UV8t4whPKmsG6FL+rN
mFUAaeNvKKySBI6o5fOkRg20WweouQYohHvrul0DeGc1JQiO0Mt8/muaDqbgvEcfFLC6EvJN2A0y
zWQMh+SDsfbbMVWSpXnL1SQcpV6HwgC0upd2TEkym2AxELv0okoyuXlrXQPpVn2LDRF/MhFciAth
9i16STi4URc0yf6V1HpZhqrTCJY0/YEJaEL2bbHJQYoOnSSRMZ+FZBFg957QVKnsmdaqqPmGMafr
kjpt9jivJguiFzwJYzJRj4ECDb8CYA3V8+VRiA7gddMlGTPiQmBhaTQt1WbKbY25unKCJWEKmuUq
3422SrKXArp1gqSEGUxH3jn/cf3YAF7nkH895rR1fZvj90Dc6rmhGtDzo+P2Vi806w1xehZAjFjX
FBqFWlahM4SNHOVvrGtUFY2p5szVq3Hp8TH2bN4XM2lFO1GAIUSpbqOI59u+UE9UvsTukV1OTH6U
Vt2uPFwR0Y7VbTjTxHJgqJN9NJOLApe0FPwPwqRfBBAjQnqNYxpPBsj0884HeHB60aSeI5umr+E5
FX+kZ8jEL10QSn/MmvsAko0knklfRyM5pqrTKFwNRBdqDIbg14AC/7V91TRLe5MfB2QKe4UzGBp5
7YXfbmeOqVCwBBvDuz3VJO1AALQ0vVv2ddxAzthi+g3GQI//ENhKr0DYkvrHqDCUzQ3YcVSr9W9P
pNAzpDhMlANJrYpnuc8463nZdRmkIDV7IdRDgCcHrpR/puXBf8NPgiFid++vbmY1PCtfKk8KNnRA
Hid9PONSZsC3uOMM+0+NIh6dOJ6hNmHr+05ITsy8/W7Wv5rXtSrI6Ohm0NcBqJGLQ6dlBe+9watx
R4AcNum3/1q/MQxq7QoObwKcIRYouSGNkYC0Xu6/o7qfDXvEXJk8NHWrYQa+LDD17OHKANM7FgSl
hXQjGuUv+EHHAFZaMkktRzkoDdC08CPVDbK6IWzTsDs2Y/6Rd0mErcmglMoniG17mnJ4yxSM4gte
ypJm718/4zKQiUi/DSbfdgmz19GPSusRhy0vIufd60K4WMqRtE+mEi/nDgcr58Yp0lacrYNhIrfn
43MKX/vEXezAWluSc6ivyrWS9ezZpAMs9+fw8WsEBuwBgOx6sOG/i4AONHHclbHZUfDXz86ae0fy
HYPx2miWHLPiBL5XyoUkUj8JL8X14XzSjEF1XuXUyQfS1IzW9CqrWNwKtuvH+B/jhXIq1pImkQHj
VIYcAagMEdTXet4QooVFF5NZQ1vb4kmNc0YULM+OR6iRdqDjkYgQX4J7w8eXW8Hm/LQLE8fvV5+n
2JZ2h21w404nBpee3mNYfWh6/oSzNoEbkydr6IGS5h3nXNSngsPDU3XF2ug8KN92BMDvQmfkhmfo
pw+tdHUzKvF2qrNpVccaBhBGC+kD2fYazdzUJN/TExcOs91XhXL1IGt15jUwL11CunxYE0t5dJjJ
9bUN2aL4vShJeqvG/mv8rbp2PNVsuC1mifTF7J0OZCSWQnLhwoi3AKHMt+5b5uLeoUhJrvVtj3Ny
vOxbR+zCrRHpqJ+oOVAImgUbzm1Gn4+Du5UIbOX4F4dvCYA5yxP+bUZc/ikAUrSzZR9Ds829NKYt
UdUoay3VqMGc1FdXkmZWD4b60xsIKpyK53gf3Pdvb2Lbo3i0vYH4br/VrnONXm3GyMEqXMJ9bBtK
YEtb2jORuiynV/85BhpUcdiUe7XXaWo+dCFEFIGBk91ax7/lfdQ3Io7VQXBczkIDdUOgzMpUxziu
saD1OkxZ7+psqqjuleha4AEVapl8dajvxkJTM7vV+msk4PA84e8Drt8zuPBFqVQ8KGzq3DSt08gg
TRu5u5rPSDx50SUeCfEsIoPyJeFzy+jxHeRQ+FMPFwquOS809gmpg+8rfB5PAYaLzNiR9IDWwKP1
QGEuu+Z3zGfth/G/Q3l1DDG15D5d8OMr9IMsGC4wMugJ8B3vszh6Zu0FvPsvrjuGou2iOX57A+8P
g/vS2CZ7tI09JPSKEcaRMzW4S6ie/OuALw9DlqGwJJQ1w+Q+prxR+44k3yKYJ4frTd20LL+1qKYP
bDGH8o12z4Nf9Dr8YnkhpQHjFEtjj5nvLj0kw/SAIjeQ+SodlnA/2iB2iNxtSvLC92CBsV7RWW3Z
zeLRY9X2l0QY2uM0o7A4hPARxXn6fsxKA9pjU5amfrzeKyx/d5i+ToSTfaQqYp6Cnmikdkx+HLys
7W+tbsX4Nr6mLaY1/F+y0MjO6Qr3HQppBC+H7l9Nhs7gyqo0YW3kXNbLnhL7EM8EUPdicKzGmyd2
VDrorhC2iX8VXpjFAVGpUfLYUz+yLluLK9H5EkM9LEQzLgpdniGN4DGxPXIieQ7y2rtxX3XIDvhC
BXSq5um5RIk2JAiom04vjxaBlUyG5kZfYQGx+wgmrIHUfopAnJE7RIdu9TQS2+dYg5qHhX0XKsQE
g8LyAXYRlDqUyv6YYW16qAaX2AKCNPrduyn76DpJfWKiLj07Bi2TK57eKViJhInQiyn7xa6qaamG
N4WvtHEvWbIcBFQUIQoKhrQW7Yao2rigSyKjlSu2zbPjuoIT+uvJ/89z6D3LtIIPRYIF5bXeUu1C
qmLe8ssqP38B+3fKDvWV/SOjiAL95aqjBtE/8BZQJEri00mwWXC/iH5PWqDPa1yomsyHXvoj/kRF
DA+REghptOd3fl/BtlX/WHTDej/eYmWF3VipSbijfg/X1+4e/F0MzHITMJ4okW31BnTy2HkbB3+W
acJN0TeV1KwhWt/wItfabI4hziAM1qR95bA1uDzMt3G1T4fFje/CcWaPS8D04WxqL79HYreLE6bh
QhWex6jLKBpfagpohuygpMP9cycauiwdJDmeaM9tFRHoZjAtIgCe/HABDmirxRpmQnDiaP3/CqR4
u94e02/Gd+WUkVfN0KlC4HARAXGCc4fGiW+0xRblGg3PFcFRQezKKfzrTZETHofLtdKU7AWXEIdt
StwUgxJmN1mbrVXdNpH51X002ywHdkJ/dxKyEJ+rtfpUk4+fwZKXGre5L2DC/HCLiEzGmUF4LGSV
tCoCwC9lqqtBWnnSJJZfFGD7jnqBV0x56e5CqvZt3dYiaWi68Lx2NQTuYURs1kRQzo0uEjSgtIZK
xQ+HXvNGdHsHe3NaAuYpkDtGTRStCFidjMKpvmiGVNuZ1iYmNOeXlRQYodTIbTfP/T+R62B5lm8l
ixQwQlA7oGyznVErLkQyIwC6/+IeuXiFb+4GFl5ZYte/+7ArYckUcuWev6jCoUFipABjGKEkFQFt
bamqNdUoTzGdw4gPOQp1reTH7KK9vb+pe7z058KbF66WyFhmaO+UoKPP99O62fIfIDMFWEK0yzhS
cZakGdEDo03CRf12QMw9e2E1LqS2TZ8LLybDRF7MDVQT4RoHCv2AeY0nGnlxFcf7JmTD8K2PrMNg
2GlsgimamDzKP/hIwHcoWEMKISFQope+3XS/fs5V77TEAkxtstmM34WGRk9lC52C0roKr5zH1ZCh
Zp3wKYRPrGXQN+75pxAt+F2y6+Y3EXa2S/UA6BjAqhWkQw3E9JwbMHCuVKkaVPap8ETI3HJKaRFj
IMUCKu6hx5qCf2xgTjTmI0G+dyWLHq0WDPSROswz4TJTx49FYftoG6kYj3C4QkoIyyYhPqVOw1VS
hCHOPXGvn99HCgPPVRBYPLRXPHZKtQ48mg1LD35zCY1KWxOM/+pWBmpTUOEpE4tvtiHf1JL9wZda
fgwofADgxaRrjBad3JvKDemfX/mI1j3m/1wBS6WvEc2rwXlGX7gCzRfkjN7PjgYJFO14SD3boHjN
plIYi+n76q86BAbxT5398gdENV/Ru0IP9ysNS2EWYOmMngTcITxiuRZGxwIRZuXPVQFn+Ei3vOjY
sbgJgv87uIQsRUEYdQ2HZenvLKARu+Nr+Nvzn1w1LScrXufglQnm6ItK0RUoKb8r+RhjV9i5fl86
EL4nq0Vkiu25+s+9bq/Nb3CVO3cZFslL5MqIOwWaGr2J/g+PT5RbVFN5IqQ4X3vilh7GOSZYZbCe
k9zXoz9diNApA9HHEgDrqnC1elN/VJhIHWFqYxhqonWEkozIN5w5qNvQHsMTL+4cn85Ku/jEHpHE
iBavzAKDGoixSC0akSP45E2VIkTpUWUXNzB+sGDbfykRF20I5GAg7QAf6luHpwx9WJC3wyQc1piv
n0PtlSMZYDvzj/XEy/LwCnHhgbmI2+314hinLJJlsU8PIcPazB/IafyERlwSw9ksMgHu0doTeO0j
8PQsXYxJF+uPmwd9jZK9DXXeu/Qmh9rall35P3HtreV3xbzAERUr1eeWkqkVcUzcgCv2NtLS/o5p
StRotDCHNxaVAebPvcgdB/eZTpr7y5G8YzZ6TfE0tkPS5mRrcJRPkMKPlDbgS8iIkTeKMaKQa19u
AXq+6rkahOeHiUdKMsqglAO3Xiq8Rz7WjVi6TZMTIznxYSq//q66E3R/jU+0KsUV5qd7bzsskil8
XxktSN/klrn6AF+wux+InLFO4Mu03iHzOMPluzi2urpq4Jkb5VYgodtWaj61L1g3bz7zRIcs2DaA
IwQU9wNmBblxAvj+3z0yeOfI8WyInW+9rc/EK7K8GJlxHLNkO6RJd0Kap1hP8yFhGaBHTCAfBrAp
qwS3z43Ao2OIYoA7oX1KqRYKWdDFs7H6as3tr3uluwsv2m9fB/hY1UM9sxuU30JG88WElNSoJB/1
mE7QptLWP+Izbinb/AOOhErsR44wheXlZbZqRRGcMzgXFP/at/+1ZFL5QNAj4V5XW155rPBSP9LZ
M3ITSV5jFCezrK54rVp2zksVgbPVmexoExsDYqUY/hiUyqFFX+xrzlm09VGOERk/7VsjRPYH7RIi
s4qQ5xryEAwGztjbBtLHNacQsu91DGuuKgZaW1Ux2344TvdOb5pjqeFhTjCgpr+mdeBEGUUCpvSf
uZDDkz3hU+prdHZsi8hU4ASj/4kELc1oBK4c72b3WEbETwDdu0uanzhQ4DYZIE9Uap//2zDTFp1Z
yBHqyfHsb6P/FOvgXDjVPJn2Sc4DK1Awjq1ONQD5XBjtshLwZ1nRMgsudNJ5LiYPzYdwOE+VzI9Z
ZPzdxLxjNNY9KzhDX2IY5/quOugV5khY+qjnwII0vnM1rOPThRHZuTYon6CSvy37EejvWbWXgMyX
b1kOVXWyJ5cWTolu+wYFgkvXAwXvr0WL1EbRpLtfv8IcniTsNdgDZ3jRScESQyAYpBHszl0k4VXa
dF8Gk/oc8bVTHzNNOhTWuYV3D5CHI7NeeFSqFSoV/j+DOjH7VziXTpQ/iU0lhJ2hNeEROocrkUGZ
KofSVWni5O9Q6/hQq4EoEvAi+wBsUbE7xAOGE49/xG08O68eQDFsSYodXi8Y3Nrr9jjDU52wgpz8
cf4UFovE0NOrX3z9q5Gv9tQk8f/Cwh8wCB3/2RayCvwXVXrfTCt1gjfOZbZwmRwM3hSVv3KijuUb
rjG///2/f142aYH3WGM9m/vPawGoMOkO7bphKBBxUh28b+7TMU+MpaEjcNhWT8WAhecvpRnxV3/S
X7E6oKEsZYUmbxU0DH38jYKyxU+cVTwYPBhXba+iB9erpA2G87y2Pb0ZNSq8IOwts7/PecoZEcmB
EwGKP+zHVGJQWC0pZHFj18U5prQXIA5/yOC/pgPTtCB6aKe9XIZaXjY+vL/0LP2FMK3cVqyf3GL5
khQ1xlzQQoxPg3yFByMM9GWTCQJ20+Nkx0yu0mklXm7L3rnOMmMgor6+Tnr8mQ+m5xcVQzVNwGaC
rNTzrbMW6wg676rpDr2OJeRmIHCV7Voza6KdBAPc7DEL9fPIHhFffxsXBQZhsgeHQjYw1qGpiO98
/fTR88Gp3iBvIpMfM+7CpHq2TWJ5YYcBAsiSRhbXsHe8SPJfG1U+pRt+S1+2FDDSj7yNDStx5MxC
0fadk53aJvbUeQNbZO/AGJQNKZ0FOzmEpmyt3k2vPJDGqbWEbhUpS6seoJRgtXii8tU3o6gYrtQ0
Bz2zg1qEI4gWwlaVJMEwUckAHArtqfCCQUJ5ZONa7BQj1lvgf7KxsxrPx7eUoD2kAdQlUcyR+T9W
keRzBnV4Gimw5vQS3XbPD2enhebr0FCSNcYsMdHE+E8rrQj3iHs8mBuQ+sVUqwn/xXBtlyAdcvMO
wa52dL/yc/jOdGGXDExk4cZq5lF6jgGvt4YVB9K00HgUiEFZi4XfrmhpdwKbMsdPBKqGX0rrtAmq
ey85sLodIIDFrIOdugDL7wY4MOfr5CFcjGIMY42hFOTRH0uzEkND+RMhfGsiOvTDXrTnvXeuR8Er
s19LsWApuQDolpQOVhy9/dOmJ4jZl6PqjK/K7vf8b2vgsWRi3DMTdKUvOeO+NL7CHFrRmIYK51kb
Sg3bVE96o/7fPXUM2wcspilnryjmyEgUwWnU+DkYl6c3Lvgut0qY26Eq2tNt+By71E8BjRL7373l
66M/rSDrnXQihLnW7UL58lYNghU0ME7PXdoPYHGGA4llQF3KV8eMScV8fYPfGjqx4XGrE1Sm/ND9
a9bWCVtSNtrw4pcsPmWzwalSbV5UVHvqwZ93BBrIrY5wXeyaBAxU99rYIyCq5AZIOTPF9vLl+f3k
zybTBISnAEbrtV7+4S8AWHULJUawiOViW8adKZN7F28tLtzoWZ73kTkT8HK8V/6hOj1lSuLuh+wj
X7PQQ9hyngH5bLtVCVPToZPP2BO3nEg46Z4/oIGQAflhLFU2yZPKz49+OkYsltbNLTksQCOl+EWS
fBXhIRnLbtEAkqKB+ymn9lPUcE+O8qzSHwEGLGHcGKJ7lXhE+xnVZAXXNmXw5aGwgYX8wBi91Pty
15Cq9JEU3pQyPZJ+SCB7dE1HG5jRQjn2KpCiB8KKmOZ1tohs85EO99pnVRMHoRmkpv42PWcXql2J
tuHe3Ix6REPiStv44/LsIdoyjxWU30jOzRJukv9Pkfw/1Or/fpinCK4NxCmIBj4X1cc2j3YKgOJv
k3/xaairIQGltKqnbSfTjYllxkIZH6BIOzWN7otimAVW67wrmiAtFBCNCrZf1U+wAQR1OBkCZw2c
TNJeZYu2wd3Y7bkZ0NScpRdOpg5blU10jm2ONm6xCv9vcj2gbwIX3tLJn4tFQ+LtURyaZmXKUVtk
DvgDLDg+RYIMnYoEItBMyW0F6++u33EYHkI/D8tVZhkXsAoxUqszm1fYH9NfsCMl42adJi9zS5Ic
Ha22c7Y1mV2drcaWhM3SU1kS+O+5ZzVRnHofs5IOqAYPlbLln8RBixY5fhozh1BFLOYytr8pb9NP
nBsHzzX7r5kwMn3imntSEGI6+gWu2CIYCIOmNL8WYABTGvx2HhS2oRZpfE06yCC7TPhtXmLyHVKQ
LKhqL0MPNtuSP3Yjptb+dUNRXkK2hQzLdnG+XyZ4i2iknXTEIiJelak8AhpFjrxpo81pcYhoc1eA
tXtfdJ6GpP1r0lW81QpOYL0XgA7Ri4X/kHqhm15TwBfXpHzw8cyfcdnm23CupoYEczWEggx27a07
oz/dXXR+lUdQN5TtnJh0OLa/AznHB9SyNFQGCJJ8On75I4SHyBIr/N78QowjVbhfQTHl+XXXs/Ow
of3qoe8LkVpB/modpBITSUyKV9gUZt2hH3gEqYCqJN/KVKJ1eLMEVxgKyIfxHAUIOlbpdSrgk1ZS
PeJXnV6A7KboKKCHuf+OWHSK2lSFILRpMmYJGP55lcFyGITkkmaldEyz4Zz1A+P1idCD5BUaM/6c
+DanDyLoF2ibbTvWwnyaaz3GD2qHxciv3WD924EAkhz3XLi+ECcQ0jcIDBA/API6u+3T9LsbzzoJ
THEplwGekaxgfmzgwBhGJkpbtfqmxaCQRmLVnF4EKsNiVlhW9e2aA6Q2FSJ6ft6P3eyzjKGzEv9m
vr/JzEPSI5uSeZkbLp4UCrWAF4bXstviW7j1QvV8iEPEcvkIEMpqKwofa/Ox186/iNVRBswGB5FB
VmB6g3Z2OD87d3fDU5TnKPZohRtSfpqeJFodPeAgbTIKvLv/ZDs/QngqkVyoRdrhd2lJpDhQ83oo
MBiyjXphkMQDs1r7URy8po6A/eRuyI8FW094gNj03CbPQbg8zPCkjpwftP1pWJile0nqBC6jgn18
wYVGwPwF66Ggyz5llJcSkEPkLGxYE1AzNNCmYXBjQOSHCdHzLVK9uvXfUCwyrKyiVQJzMky3ucsh
sH0V3n5a29w3OYnFu11lj6i5wvqLPJUWUtI5GJ4BsgUoWd/F0zmG6cVkiyBftsibui5C+B0ypp+S
lfWLvXjCr3sDlSCtawYZJCt2wiEzSTBoEOnN1vH/eCEiGrE0iOEWrzxO+sQLv1o1exex4qRV0XOZ
uMMDji5dR0pazxWHBiDajzJ69ffJvaZ8iOprj18C+ou1+exo6cgAjynzRgBgyBZ2Sz41aa94SR1U
4XHrgwW2gHC3GJvZF7Qfs/00NPl+BxlT3P2kea78jjAC9bQGXh9stmCASZDx/0TuQlTZiSx0U9k8
MAAhX+0gyys5mCbxYx5Ekvf4tD17wsW/oORjIVk8pBLiIY5nALChgn6xjStPH/Kis3wmphtkDS/9
6rk8qQcQNfg290WWfHbWXWDlMDvQG3O2E/AMsdXDuAzM5UAzYzUNoh1YCtZp8A3P5VSAE2Wfa0lQ
gkpIoZbjRgbmppi+mcp4Mua/InsSLeBi8B/xBCYE+prBZ+sRsdGT3J2RlQxruIQf0Q0Ft4DC2P58
dHhfk6zD7oVhCzmp9Ze1vJfW1n7TXIDOytsLCp4NTDKvTHKPoz7MSravTjvvpWvDNyRNhTaW9Ohj
0qCJ0dRvl+6o8UFQH7gKTvM+3WWyj+exUXNHMyxGKm0SOMqf4xMkwz2auMU0KoWZ1sq9eUYKQJ9M
8szZkr7s/6teuoO8ZUye/MvkQy4Wi6nU6hpj9W04LApwt+Ua4J4NxwhgpI7WBwolhCeNJVzrWr+h
8NMS+gg8b3/2m8RnL0kZ0WYCp39Hj4lkTzFWnGUSUBSlvWFNw7VHTWpLWnSe7izNi3OUbvRVvb8O
NzPQOANcEFUT7mM7Y1H/F36Az+OjJy5buGtAmGCVyhW53pITf2w/fgGGtdzHRYE1X1IQ3ULuD2lJ
naBoTMTJXIGeYSv8yVFSPzvhCWdYvHtrDs0PQduLonpJBw65t89881hU+CYOAbZTh6AIHIr4YwG7
TTe13yuUvO663Em1E79yV7cN1E7DhmQcoatImTZlumKWu7joAESWKG+/UyE9x36sbgQjHZaRvEXz
MJqQkEjp4eY4gHDro8oKTyZO0lU99ADNp1PSd9hEnZBUROxJsfrYvE1C0WipiD9vIFun0joSK5Cs
BNHw7++gLAzo7WfNr9AljCgOQZuBEXQxyweykqznmbHOgKVMKhnhEe1FIx2x+H9x5uF4ah8/wYf0
rbw3sGKnAgGLvjop5M84lJsjA1FCtXkgKO4wKuJIU9Y5fZdKGSh8SJGzt4FGGXG4/HkW88Gkfzuw
OykWY5DRhaLVI32Hvjk3fxSUEX+MQmoo5izVh/qoxm+9JWgFKNz4ggCuwI1jJFW8QhGq1pgggZnc
Kfu5ILfCOj93p80ZC0PD6S6wq3N5kGQ4QGR7LVjRr1RPLRqsuhbNltECPGHWvtoz/WaJbBPA+B+n
NJul+iu1TXCsrIkV4r8Rq+4UNFd3G93dg2eVTtZgYWq3rpQ2055RongFFxCux2Nz2OqWjWJty5C/
PIdtGQBWgYC56v0BJi+gJaCZzA/HIAe33LvvNO9MjMAH5lXwZGTR8t81FfYdq9q/fqGhqjwUL99N
/+HdydrZdLSs4Em1n2roQTcBZr4L9ZPwxILhEYoqq6RU2HuHCkqPTqtEhz4wmyhJqV7wmOsgeT6s
rFYW0rYbRrmSg16Cyvypl4KXoKLZiHs3YdDT7u1ixt9rrt+NXewlTLsJBw+vu3l5pLdqCmWPDFUs
7xyLzxVo7Cu6CyXgaG9f9V0hTUqW/GC3UGn9vDRr2Jv3lG02TJmfXpye4vQt7pW/QT1hE4VMwdIW
0qS8Cycp7o6knf8bnU2Oynp6JQP7qSzTQmGfQXquVfjL5cPFjhVxcXbnMczM6IkXxJUQa9dzzEFp
hQl8wT87wXjIiGcSYLPv7zZu3UjOWe7K7rbD+x8W0WstecnUabEXVYQjt4CKKIXmnOKtO+3irY37
HQtRJCyJCiGbsvplJL6oJrqJcJj9oVk/qcLKivszYfna9j+9DGFVNw0VKpewYXtwW7K79SCH61KO
YtietPgUftxJdBelkrDVCQyD6m548xs+1d9gmvto3nsX2ayLuVsKvWiSXta4jdYqPys6CucRpolV
QB79yEw+M415kWIRkMoKPBjkYMsnYvlJvLG4cwD91Fv5TZ/R4eCGWx0YZTenkcZxAYiYo0MlfmUp
3vFLCKE+33i11kQ9RXpFeejssQyf54tngRKHffxpR3ALnyzn6VAcBWdkrF4BA62x9MPihvOH2YHM
pzIrD+nzWgKR6iNNC53rUQvzxRdQ3jJvD3gQ9SeDUrIrWtuOEY4yVWCWVJpDPstelnET2pHJarUb
1PtVFx3OOPsF0I4Tzo8wrwahb9NTL9aphWgRWU1JFtDYExKn6i7+TpPsrmIf+4nEEcMooWpk+RuB
6AxjJaxgr5GLCDmCGUo1KAX0+KjnN4BiSWLAyZ+UcpAMPoiaA/z4H6ngNLJduQgPtBYK7WU5XLU4
yWxGjjk3+jV+9IPcpe06c8fFBJGj7vFdEvvT4JDfu2gs7fXMUqMNuXdddK9wmMXm+apYJKTpoSg4
BW+m76WCoPBVpFM5DCXtY+/PoXxf81LcMY6/8Am4MvLyGUzhyf7dSxvYBaL/CECAOQBn6SWzFWiz
lbUXrP5OBccVL4yisgrgKMzOe8O70jseBs0ZyibTagHioyvoUO1kfLm7wmmBj5Fr+HtoNSBde+82
IpZOS7kHLC23+iIFK7LfKVrn8bwAYhtQt8K/RNWevwmtVBj9DWSYfGeFwJd0i8tU2eZtC5Ypb326
7UWEj24HSlHHQ2doHhmOgPL4dMFh2q3cahIaOE+aDYs+zwkJK0BFjmBpMnEm/7qnc8A60S1mivQu
XGZKzSYUpT3WZEDmSue1N4o9y1GNBZeMA44m5uhy/BK59ZdIDxivy+n/GgvMo/mHJDE2pex/i2JF
Ul6NY3r63MWl5tNW1b3z9Ag33C8kkHEzwOJl+adYTAQhQLe9owiLUBPjz04izbeWC/M3G7x7Hri6
5cYWWTz4ExV+Bsb+b5NhRO00yapJhB/9dQsiqAGs8KumwxOqfbjthZTfFoDJS3av2ktSTjzNyPAA
mZ0KZAj2Kazn+CEo63pyASOVBD8frxgT7+vlP4LVhGUOV5GRNAOxwuZ5fxoXF+0/VwFpAZjlbEI0
jbnwkF3SpN07zpQ4I0NH6Oznqr71FRahAhnR/ghOMtg5T18Iam54pVAXbB1PIGlBacPTM/bi16hV
LGaweqj6B1aCmJB6gf+piS6TULWHhgOsrCpitqcIng5ADhNBA29C3J0GYs9nelN1ekTcR5dE+LVi
F7/bXB3oQuPDQZzj5yajuzJjSF5JaY8pB4Wk0ca8hMs5LT90YIZ5Ovn+EydIyw0uz4NC+NRsDB+I
QXpD6PUV5O28qg1jr6Er6GQTnnl4xp3EEJuqIafyEY9U8MzjrYQ2Zaj1oGkfJYnQwkPxLNiJjag/
WZdoxTAgKSDmhClYK3sIQuWxBgB8K73IKLM0+ovywE+PtNaVMrlUVqAJS360YWdq2bv8RgBomJrd
lvXzQWhQeLUvtCAhOBlR54tTNlOLop4FBNyRDw99jJMT091bb0IktHRh+52s1a36qzc5lpdcTkWh
hN0iywxdc/hus6fPDmlRcUrjPcYnILJ/Di35S598MdSW3lnzNZ5aw8kyrlipSuD2ZUXfPfwTZrRz
PpO7YQtOBQCraCuaQP6074yfM6ZoML5QOrAPDadPFztNl+LrbY2pWkYpj56Rjo2n2fnU0VKd6EBA
cpTzInqhMwLgMJP+taHLhm3EX41QQ77cbDSIE9itFNtjUn5tZSrwjzovQS6/H/BKGhrVNzvwPBcs
WojMcN9+Gud5ANJB1GKhfiMMatHiUpwgFrVijvRpZ0kti18Pr6CdFWJ8LPIvUdIzUqvnI31Iku9f
cKQ/tPufv81eqJRTv+PQSXcl9Jts5qViR/3z24updEuL8DB+IpEOL8Ei3x/Nh0ftBI/4ypSIoJW9
MN1Gql7IfeAU3tf0nRfyHjxms4mjckV2dVQwG7hdZk8Kh7IKwYhuaAycBz1GbeYv0fw3jd9iok2p
JKMCe4e1gwsHBebYmGYa+KMgRqxxl+vCk4Wh3XpIistj5XiGQQaL4dwHWG6cGeQVlZo2LL/jCtlL
YcvwLd5H7XglCYzyL9xybDjeQ7LU+wi6UNBg4f1kbeSt3RQxH8X9ytQUrWbYerpdcA/iKLlLEjPa
gnTiFoDdCQeyVi/yTG7oZpteB1LAzg8AkbmbXu0SHjrt8mt4wTrxNqSqz4vEgZ/jlfX+rUwirMlt
g/SzQPAM0rHn/d2t2jMqspg/VBnmm3LTkzBZMu1H1eJ1WDbHHH0r4g7KdAbqt6Bu+97WAhS4rusr
EfTBDTL9UgoRyb+39HGNWjGRhee15JZ3ss11RTShQ8WePNyYkJIcn2J4ZvMfR9wR2rRw6sl/P20u
QBZuffHnkceAPYFCA2IqI93MhsoX5RBEfLkONFOPXtlcULgeFzQPPIKslKL0LYbLhZphedz2O9/s
NoXQa+YQMTEmyNoSHQ9M7W1l/WsHRPWCRvz1Bi96PwzJmIwOnXWqKUfDf25Ie9F8vPFB/a/TaoNN
OozEW3Kk2XGMns19u+sWeM//6sjkfzx5y59y9ae+lkz4NgcO6LkPeVWdAnqGKF0IDjoTf0nF9zcs
a0ybLAbkMcm8Qtcd3SjIxsNIZ+g1LqE3aJxjvpPTuSdlZ5VruGOjHaE+7EUIw/Mqx+4B1/eih1ue
+Pv48OBjrqX3gqNmlyi/SQOc5488nstjWNerxFjYabfNB72KbiHo2VTPuTCXMpp64nkU47+ySZP3
mlta9cfzRxX3Cdy4AJgWORRfszG7PwyG+AGJd5fIETNMGobTXT2WbgLh37gxhwUo7pTXZvL7cym8
j78S7lOG2/FmIePwsHY7+TDAYfWh76WmVhzTBi/vEemERUTLfU6ZfvkOTvfORBD47xgILYhqb4kN
F/wNeu/J2z/tDGZhKeFlUvs8mGEGzXAyRXEY8FTKmiSknDOxLg9ZUXoqtjgteLnok/mWa/tnHUQR
BcNwi4OZ20F9HmOmQdmTtyhfOtNGlV4E8PoSQ3QuIF02Rva9zUrgeX1VvYrt5dhfmXdSaiehT0Qk
cgVvsNPO2svKHJFGwvJkEEw24hwYdTLui/mI5rBC5vDZZ8Nus1i8KReYCVCudpHRMsgZlD3Es9jt
4Sn4t27KQJakLOufajBHRAxHCuf7rDDmhl6SzkJDxaAiAQmvNBCTw5b7XQ3S7aLfrVLLI4Ny8YSn
ZtgnBUvCshGNHFE31THxob+sVCkNtqW7S34/zoYYcWpbOSqb1k3OcI6nYm3hrJaNHKYD+N1txYwv
LWncP34ufap5VfBYxr0+v8Dk0GbLtrgKKwHhhiasKFgNjNZp52R5AXnRdePt0bl1YW4pshGUcDRO
ZOwl9XojdcziAuCq/e0bpJ9XlF8SL/Sh1XKOn9U2+BQ95SBVhE9/OufcBonTvkVEwpbRdhbfLozS
5IMmf2vCa+a345lc2fT6jR23F5NE+g3zLQhG24CoWy+IGZQ7Hu5PwgASxoqE13IPE9x2ZoDJWCZm
B0afNKO3aFCFQQtLox0rZ+tWlJUq76d5ERc9PJxXPS3luoSDZgPGFft6x8164efQ/q3Xj8nZPI+h
DXIzp4vuxYZvksVkEpo7qJNxt340Ve07sZo2JJO1upvqZfHHZQFFZ6Xk3x4vk2AS/Wr5PgFIMesT
J+cIF7EIlk78Lyh8/WWwYBDlUMoyIMR4nC6oHI+WPvjK9OSXGEdikHB92aE6HgKewUvSpkZ5oCnN
B69JgW4oG2CsaL5G/CR/2QIFCB74O6ADdVPnTuhKyFCV2V+8Ld/sB5eLqtGdEoRC5O2lc0xOAlcM
c3oh7NsgMQEUI0TNsVHg+/r/h3i/dbvFWZkJjjhkU6auwSJX2zV9BWcQzvR7Qv6Bj2mVA0TZkeVy
p3ewCQERbzgk23tTwCPY+8NWQI9YPWFlethXrKj6r8ob2xG+CrwnNN+Hb3XgpzKCp5sy+6Jl8Ivu
1QxLnOf4+T7/cFKdRXxQiv+QEjExWfbNvyoZA3D+Qlb7QD0eUsgT4uZlptsBOKWYG254c0khuVFK
0A4k5rTrTKoogfu0y4tNVXohReI37CxW0SyRAx6EulpFXTrOHwUTlJjm/fJPwnur4Wc23OFv0d1O
3k5+srW+Z9wV8snEbhwfl1oIxIr05TsewFJTRM2qWxMTzoaVBfaQhe9eW8GVCyr4ivlgSeTtBYjC
zOPYOcYzsHOW0QXOoXw3xx8Z+36jth3uPLAU2QxwQs1p6SfWMCqj3hS7OqAVzNQd3R/RO6QaLeo1
5XA6qKsMwaS3Nabym+QUwo4fT4WrbU40Zi5kWoROCBlqqHbuUTJOYE54yzuYGIbz6z3lhSISdaHp
Ww/n3AKBTyqJngDbRoa3Wy+cthirIZtp7fx7HbJtT57rHi/HwZquXh2dczSUnH2w3m5CrZHeUG7S
dNnwHgaq1Czoc6S7y86uAtSGih7T8XCKIyKZo280Y6EC2PWtsj2VvrhnwnjvVsvQU4VIpRIdXkSE
Dny4SzF1sCan3S2K4xBZXClzLX2gxyzm15tDfVxu4DMV7JhkV0YD03v7x/b9o1i4m8W2Ca2gdNOU
AGnxJNhw2F6sQxGlm/1j9IOhEzW/ccEWNfH3RdXM4nqx262XS3Mdm23N5ih4FV3cdig+q/Wn468G
Xw3NcWNReOD3PFsQK5+NVxLEVpkg3quGcc6PyxOoIGQHwpLkAiN0zV2pNTaWMvHApjKEngEN4eXQ
bETn1d3GWtofzVHDXbDulUU1tV+nxOMVi94l731L3QNo3HICQwbHgqUt/T5OwSliQGk+bsab6UCy
eb3NbgVtT+1cKGZ0/hwkaZtVgad1MWjzg+5J3ENfihmgtuPwHipOeS0N/vvBXqYGoSncx74IPv/m
UGYbWkD1HKCo3XbcDJYn7+SLw3IoKbykRD7EiKyqr3B7phjtgBtB3rd4xLOtALiwiFbdTRlkf1Th
8hH5/XtkXtlH9A6rr9p9cSiNv6Hq1PvWKGfoCroEy9zkL0eZPa2a3+H5TnfwlFAUPWJj1hWH7a37
HejpPKhM6IUpp9NANgVTLbjUhMezlwUuIqNNeLWgkes5RDosfeuD8lvh2M1VamWp8QlHIBazTors
iOPCKIkllZO43d5CH2Nc3Z0PRcrWF9C5YzpE9jQoHlygZo4uZeljjMUToJP+RXUnah9XEVSnLwzp
E87n6dgzOukofkzYHRC8XNMlv6W5VHXwufnZ1vK+w0+UNC4u8x1VdZoFQR7wTfNsfHzc2bkK+Tye
JejO5QAi+Pgexw4y/8ZbID/C+7BQPjsSpYChRdwae/XAwPmDy71B23mzYN2Hi8BFSVrPIheIjEbx
zrKNMw62dcEyuDCIh8DzXsFE3hkLX+uFhXHnjh2Tzxa9l1pKsQ6U0/e2F6L6JOCvjB+O9i8oUtFy
GWPQRxAoV4n98QG+VaovoLZdReKr3y1bchE/Yy699Cf1Gyivc6EruiSJeuS7fW7Kc/PFArOhwMO5
l0wmp3WhSY6n6maymdYQ6m+GHomE5gaZlUIA6/d6IrLC+J/mDIGMYd6VhQoF7dwpKT3VgyoCWfFA
eq1iDw7oAZ76PSP8S9FVA9QkHhZOkNvXDmiJEHXHwWU7g2AtEYTY7fzyWHLTUjqwEk8BFEvU29Go
8zR7w+rnykpLf8wT/16uSelRJRwfepSdb/HwVr+73W8reKfU5dl1sPtpGkRtE941wCPyoh3erDkA
3KF7cG34SA0AQ1y8pFAb2ypnNrAsCvhXRTlaOJO6+2Gho+T94uKNsAOKqBsxSPHIjYzY0TuDa19S
hRzUkhWrF2JdSO+Xc1y4uf2aMFpYDhlUO9T4aYpJ6pyjaf+vaotvNQSCFiFVKhbVXc/W0hD2bnxz
tewWGvaaSSMmBsgUuCmsl8SgiQUUwIuTCljcl4bo9n4SHBEoMsvcUhA4fNj21Tg3IT4YyjX5rUbw
x/nElqTS5Iqf+yC8w7f3b03xH/l9wGpm9wlk8f/6F3FEWPRInFj0SNM0UwdVR1KxlwVKg5ZdGD+i
VQG7czOyVzUw2reOwLhwqdrai85W0R9UcJxSDr9W0Murj91serrrcEgzgkVD8BBUXe5VqClByOOz
gmr6MIKK6VrxgKzJtjZl+H1mDdBBPV/zu2rH1lmCZQi0LwAQhqawWgbQBQyn4F8z6jCNxicaXlVq
SF+C70t7+Sbq+IM8M+7G2F8rw3brkwRujWMJfDHR9T6yC0kKuNEgrlE/R9uYpvY+xcbz9UI14weI
mzkI4n2m/73fTS7xDd2xhzMvbI+yFCFX5aKElqSCWsJgzfOfYgBh1646Gx1llXR0swJe6+jzfEzl
LcZn0HV/McRkANFt9rkRgfUem7J8msTKcmiVziZzRjJmO2puut4zBixB9ib8LFcqwOaAoPCpgI1e
RJi6h+ugU66b+rSNZGiP0xVtcr3UsSPjAeMbBTQOZ7Kmxs/oLARRmz5R9NE+mT1v1T+X+4gmVmvT
gemEHNRvFVUy6o4Fl0rMDWyizSNV2pOO0yRLSLyhyHzs9txFD69lgLJ1qlcHYywxx94xroiwWbEd
DwsVkvZCRJbX6J5FKGxj94ttghjE5GJ4N6ep28+5AXYURVoBs6d5Uak4DkgLDShjYRhSPTRIsI7F
gnL62LInBrY5rK3i/3yjvsNtc8443iguObjigudERm0XjJZQeHaPi3oHipeGHfS/wIBrfne8tFk7
Xc+9ic+2iz/Ofd1kVadjwCARiHdccJpeHE/0BfGdroBRUeyOwpeN46hR31Ggbqe9TUhiXOm0BEhk
BzDr1jTHm9F3PjOQFvWIeANBq/SrTQd9aVBnVYbNCVt2NgzGQWH9+YeVjke3IW8KXihyq+CJ6S06
cpCQ0rR+C6oe4nkrzu/xXCeT2WuRCS+jogHKbkjh8p1jbtUp+vTeh9yVM/Wp1BQ+WYcPCcwpszAv
ZWwPD2VljR6W6xLwpuzNAzCpSoUjnirEZZOxSrPIYA4boN6zeeZ0vHCl4ly4N0FrsCco2udyO4cN
SijBa/VuTM2tiNUEAwWnltreraaKFuYLpvTNYIyhwYcGtOtyP0kd2MJKt7/mzNIoWbt13FS3wQeh
fqkR/Fmf45X1eFSnhfgIhFx5HO7Kij2p5Ge0pEgxTd9nxyCuYe++ET/GWXBqdW7Sm3wwGjQWixRN
0JaECGDTHmPQH6isFTndU9xO3i8pj04W7yxISlhfdElfvR8GM4Tuul2N+8ZOx6jZwNdiJlV4YcYi
zTfLnfEU4MJ+ccvCm65ltwILj09dO1jC2lPnQae9dM0GGFb3Sf0dq96fpee6NzBGHVU1L91en1gN
YTswb5pTSsHgI5ZMuh+NqW62qaLj9vxG4qvm2A53xidkbjFnRdXH8wYB62DO0NLCOK/t1HExV6Ku
j/SrBaUkP1XFAciFnSFm3uiNq3YOpYNBkS2CQrni5Pbj2vHzZEezNI1g/o4+TSM0DsiPMG708vhj
eKqmP4JGGGg+pAfa5VTfiOyURaJyuAJuHNzxNwH9Fuhzt6WGd1YRMuCoacLnGyxOqr9kFnAEbQWZ
VTnu7m56LvfkhgeES2kYvvCpc/vhgsdD8Q+LH8zScxPWpVAXRU6cb8QewK0wp0/vcsI1YmOSf6F4
8Wh/4CqP46KdNBr4NUdrDpR5j8E10Ydw/dZ9swiNTqswLa6HTrXQU38Ev46T8ifbpbS/nSdkHSIj
UMwRj/ZcFNcwQSJ10btR0Bm7Xx2AwfJRJPjjIB1BpbukVxvkA3W0ClIlKzN6PzU7gHj89RCg8Gyk
SMToOJ9HsiFUw27iZulbA/So+bk+qNrk4PjoHEcsov9+M1H8ILzNwzPgl+U6eXiyQTUW2GTH2Jzx
9cCrKAmjKb15/pmMu730A8NKA4T7Cz02Oe2Bw5Yw+pAnaBMbYuPYDMHrvK0oGV33o9qR9scNuR7F
bjJiSaSU1k8fQ2z5ep3OQf8v5Yq8dbHXf9+q3ZZR/9/+S9SPsjBERWgqEFrCEd8bmZayHmCar1rb
KayKeKJ8fWvWuoJmGFi2644bC3aPCKodJiGK2wRia2aCybhbt18/tCSNUfjBreO8aq6EM4SP2C0o
zBddy2k4cZye9GCbLtTuY6c5i38Y6drAXAZPcTwX5XWFAAIO05LY8+yD/gSxwO3EY0eg5BFE3iG2
aruDpcwM7eIB+KExZl+Mm0gbSgWFDkGsYP9KNRKj1oMpO3if6USxRSXUt4xEFYsiszo/tfUboB6v
Xlf0gZKiHE/BIrvKLUBNEwy6AN+Mu9DmY+aaPldElCaygAddJet+4VF8DEOa/CoVtwpktVlYDu6z
d+H4Pmu0WuANUSUvK533KXMdEhxUpElnzovS0WHfkHhA5WUft1XU17Bmp1nBsnRyCHocF/R8sB/Y
LN5qj779NIH6mmoEdLHADC8ER8j26CBNBwsKrlAFByDVlh7MxH6fATCXrTVcQfEueUVTfR5vfzf/
MwPg5ihgqGsx0rxy9Jbm+eD/VAKY7zj/CYma2a8pLrj4HNbyvkElKUlLjnbEaHBTeOkP9wcO4VvW
CALGFBJe5rjB/aQeOP4hP+yfVE3c2T1myGiI2Yo8IZ9+48pZrMODc/TZwoZMTxIYyrTPUKL+ydQr
3tdzb6+bZrsc+39x+g58jB1wYGo3gcjIPUzETmvYw4wGRrs3+zPf6NghzQkPFQ97B7+Cf89csFeX
JPgf4yp3TI+xZa2a5dXScP9XlI2OlwzZVOcOPz4J+bHtmSUPJ2TQddbhXccm3Ys6jOal1UUa88rn
9UVnK6Kx81+dCXW1oXAoniylF26wJUBUTKb/yZ77B0u/4EPM61YC8IIxxm+IA+ygNYCTkPEgHcKX
YahZ/bpu7KQpT5/MzXPjONeAd2NexcVTi3GmRczyUj4Sluqak4eiU0zglKVEEk+/JHDzyBQYX/2t
Iv2cVS3iZjQ+vz3hM5zcIptDsifNu2l5xFGeDEXpN7zhPiz39fB3tv5jDW9aQqy+UILx8P08naGU
tjMVTJoMF8R/bY4kw2BuZroJ/qGeJAWob5kCk1a/5k9JRyCovZXrHdNj/vQk4dEwHNEr47jD7c/Y
S+Q7FdHC9c1GxCMWcvoy1Vr0IwKKwUYhTjF8nRmaLh9CAU4HJfF/8ZpuMqiGS8pMetbJJLQNnDXO
yBNxPYd/3WWXd9xRViswYEu6Fm9V9+v6AqX5pFfWmVuQVBbtpf97x3pCPs9LaujFgZ37ogxqLbCG
KJKzBIeRBJAPDFCCA9NuXDF3lOTrlCkt0ppyyECfJEd2C5rnghm9n70yCtpMNbFAMujBnf4C6nZL
jIcFhvO8jTpT7ngwO41JLJWyFKA/1AW7afHjSyZPrEZ2ehf2Nc/oxPJiadlEuTknF362CVsVp1Ed
rzIHeP0e2BpUSG0EAFVkAnn85pMn24urw8Of3bqXyrbZfWkjtY6eDMvUhw2DtupL4+yIXOlMHZTy
gfGFZQ4pWj5s9xDqIUqgm2M7EvKgUvcgOfcnv7Jir+Udn3qWAem3DmqW3g0FR5omzZnPKdd6Usd3
2uCvaRhbaIo8sc8i/pBSFpHesa4opyidlfJ/G6Dtt+FkkhbPV/xOOqrs88WDprqTaaLWmkHwoHdI
zVe0vW/UDF4PxWLv4ZNBzQPwuEa5CDTnjm5qHsY2Q7OKQK6KNiEGhA2vS1WFnLZ6RzyBXkX9rVVZ
9RhZ07pKzX/jX80GfiD8RUOxcysxT6DIP8SFsHlxh/IfPz8kTsNG0aSsixdaUE6psBmryNlNH2ht
aMzXgaR/Mzex+KTVFvc6p66hG75sYRaWK6/bogMk82t1VBCl+8RCG8C2p7jaQuKplHiIeQC945HA
tpoiG3pGT0xXYXSdDLAu4i6TKu+dMr7GHCTj8oPIB52hjDC942Hq4mYYOS+XbG16mtc7pdkYOT/C
MksxzZh2KdrHYasOLGDq5JhfjpiANpLC2dSBxvDef50uiQZwo1xa9uTmkCB4SMMeWxCPgfOjLtrj
2mfoIvsVr6UgIQ7fcuUTuXMgAtp8BDgLyUpUNCG6KaGdbBmwjYKNfxTUqakOi10BvNzFwG2IBVC5
q15zpxi2LFWixCNxxF7iTqJZljr2/OTce7cmKBLaSROsJhow9XyPtn58n9rv4L6t+oDE59ZQn1nI
4t+TAF7r0xboSjeDV8ty/rb5Ht7hVraazWxJGqPg8UbVLLo3qN9KeXKZe4Rp9beZteAfobVkqKjZ
IT2hALUjbGiWROrPV6VveRc3bbe6GNAK2oAMZv8tQxr3EJhUJJTnHr6KiCfcIXXia2ZdI30qj70B
05QkpAXK8UXvgNomIY7vfwDJnnTN53yuVyRW6VL1cOD5N+fGrVPT0qFSVFSIYSIDD2C+JJKBZfH1
hB1fifyaRGmtdx2kCNsFBOv6QOcXiMN3bkS3dWpAPmbv/XoDkn/uBvYGO4BIOkvTQ134lG8iFKcx
tD6m9qb5keNgieZG+WcCVIceQjbnpoiU7kcRnJn/R2RwWCAm8reaH3MzmoseHtByZO1Raokbi0tS
91j587ufSJ7duh+5Kcd9kvr+lF+rM3qUxcaAXPnuGdja3PhhTe/RRYc6fTlYJdobOU4kxW52sJLq
jBmAzajn6s66nL8yXi7PfOmJt1njQSI6wVLQQyTzJssVtZhkUQre9b1nGQu+eseAgVOZRbPwwoBj
MDohvcVWC408VZ7mmMXCQucqHL+YcOKYHsmc2lp1Q6zXmc7EnWKHGc8W+aEuHRlVyMR1XHL4aULp
xnceSIhP24eWmQBIPPGR0ddYYG2NpPBqpd+L0M5oJtFSiY/Uwji2hn6vEe2FnUTwF4oni0lH0AMO
ZZ0Nt6sgJ3AXz9h2Qwh3hdPNy+rSUASMELUPFs/b6e918X95Z7zod1Uznm7RKo9RUrWbQabtwxnr
sXQUh7HRYTcNompjL45GQbErcq+F8AoilE5w0K8bCl3BKBfc9qadRN60g9B4UyXw5kzoWvMa6lSc
oeAXZP3z3Q53uFGvgsTquKWeriD18hjSTLOJGo+YvcY9lqmcNefAeRu2qqHdaypT2Xt8lqpVx71Z
P28WmRrm2ZPmxaiUZy+BCm84R51Z3WazipApWLh2lSxG5mMeGyLKnjyocvlhZAD7iOUCxLSWbO1c
2erTPtRBKnhS//YyAhn6Z6lN+9dvcQW/Lhmx+VvUJSZ6wbWbSEKZWDj7IQAHWmxk/7Ai8vAf17D1
Fbbt3sCa0r9woUm0bMVmEM+uiF7GXBt4l9FtjILDNqGczJOQHF+XsyIc3UFTthRDHZgdzqRvQTRF
gARb7n+BthHFGBzk0e8/T5Y7cvTCZNjgf9sLM6k7Dpc5Cx+jOZ7ePxocClm9P2QlZ1C50mO86tSo
05tlR5HJxW1D2tFkrBFGb66DEtvXp+xv9+NCtPRRx2djr8XrUpDpRXGPhmb3E3Gv+t/jYfvgUCj/
t2eVHnNNEi4xFKt1r0BuSb6i9ISZ40bbMjua0ZQmz4xrXxIcsr0UU9LBlm715tHG7b5VsG1WqIor
0uJPjXk2vZlA382fRAEIytkhYAhLHX8ZhhMtaZAuJG0aaD/x8iWXuxZL+VVuvZZpEh1N+9YvXSFr
vdswLyyOief6j5RbQbZlyllywvhAYsA9+QiGTstu+ynIaczPwnuA+LTYbrPDDutfioSppbx15LZ1
is2q+2OIQA6PwB9OfDrFX19RWA63BbBCpH60ewxIDRXTpzPICYpGc8sm0/7ck+ra3sEb+kmHZ14F
Y9ZESqlGjw3tFFTH1kJ5yG8GI8hbul5z98Is+1xSq1ZWr4nSMnFeaZtN05ByjLNU7Q9Dg82tm14z
u4oZpkhK1D+a0ediYZmCmLQ7inxYVysCKnrCN3oz72xmaEX9jM5MysZ3wDSnW28iDeJlCa8vbxUk
bGMATaJCPr9oD2js1h8ji7US2dQmgQldiIgSAKH+PIJhSGO+0izlHBWFb5aUGW7B+MZPDT5Uewhu
J6SbOh1BxEBBl9nD03mZx1MoSlLhchYFmv8ZIP0h6FHvAjmeTsmSatl42XpEMkmg7NjaDD3Hhd17
OIq2NF/pP9ljOpxC0OVxWiV8+aI0m73fCZsGEkeGLXKyMbJDOAkaQDUU5xhEYwka643AKVZeNxOn
lzGexg9FC6tcKnp/cN65QUmY7+/jn+Nh5KL7OpXBpwh1VdtMUI9avKAg6LW5Rkit69FV8ba0WgjH
ymvjsu3gyIaNldxjiWq4CTwo9jRW8/JMtCzF5Ktvwx+g7wJi44J1V4cgrJsH/72Yf5Aa23i8EEHy
/8XCfnHXwaj9IWxClGWnbLo/BWCLOhD2wzFH9B7xqaR59J5jC3AzlKIoaXYeJbtPGJ8fOjIEwj2y
41NSq8SjHHtTftEJcKD2tBEwQReCpAhzTyreDolaeL1oKWl5EsKxr13beyhN6mRd5H8xrjb4VoB+
1kuvzfPCPh9b/uclq1WzvLIEPgXCO9etomKx8jFpi0Sv6mtD7iG+h0fIY1TUgtx5+pFYFRwdow3l
ir+A+Yh4TUSRZ2lKKiKo9MnYMYhDuAEYqg29Fo1f+hnaRWJDx8s817P5rKKmQnbWQEa9HE6nqKDK
d5VwuiGfIJ2Ne/CsbxQm2rgPJHgUoFLQFT69228EbWxfosDC1Eo8Ho55T0nGL8aJGaIjPM6plYbW
E8KSkcL/v1fiuul502Tunj45g2o2DCy32lb7zvIN/oE0/CfONswbB61BTPvFOQZHvZ9Dj66n5ZsI
iytDwKWWWIcEBoW/yswlsvEcZvOqgHsEjo0few61PUhPzWhdqqkB5mPCyFM0reDPvwCuA6l/e1ar
GLycPAkLm4UygHQAfHw+QzrK8fHUOKJy0Zp5FWC3H4aKZSx3MVTDTDyKoXK+XZjzJhAcDwyr6kgF
6XLTpZOKLS2IYA2N8scim9e/3oKNgNQCTzFysT8CFKNMuIGb8CJBjNHmg13i5EXk7WM4RERgzmi/
De4VEMrrXzO7CoGnEMXN9RaDzhhqfy/s1AfN1Yb5qCQBa624WNb38PDj1GQbbV0la8GlhnXQo75X
Xg5PHgiQNbzJD7IN5op8KSMJP7DZJcMElMaTmeLXlE3HXQHR3FWbSS9e+uThA/hvz9GAzNycTRhx
tkQdgIE9RF1ateBlZpdOEiPROVuoU7BFvvnjkcT3Nsm6Gvwc6eT/Rm715h3gF7wmb2yThYgntwTd
GX7wUa/6QUlvaMTWVDiNQbIS4dI62Mt8vRxRIRyU3F8mRAFuPCZtMa5wxctNwbFx8caxkobk4utF
Xh1Y1xMCj1hrW7kjeNQ4Wp0FhSKSyuTz0hr9Mw0KW4oChjJFwHJp/pRpY3iqlRltQwT038KNE8Lp
dGvgcu/MNAHRQgjVE9hbJRZRdJwZhF0GxJYBG4fn9P6AdR9XW+0ySvy5Th5uoxFKrJoQU6VmeY9T
ImjiEqtsil2fhIjpFhOxwPk0MLl/3WrhGlDbAfFI3qKnEBQ1KK7lZ/OImRGTG/TeFSvTFMvUbYjM
Ac8BUOWLz9NbjQz4QuhshwqqJsvlLywr6fsb0JT585/KhdgGeOVWXGpMNUf+6hahrDeXLtejGota
N0oam4dxyA+aG3SZL8l6l/8Ykecnz1BKR++K8h7uLWsgv02kFkwYrOpR5hiruUMba0RnDl8oq9CS
eKoCsUq02sehIz6ytzPO7zHtzlF72UUdRkgRdt6PKbUA+fafqB13YXRuaDFb94Z4a3//FYVabSyN
+PXAQuj36QT9Q9Hu0yGm8SbYLhis5Te1JFafSLa/3dt6SXYXi5lc6TmWe4bSeK0Sloi6XYQzu5Q+
LRpl3LeLGVU95d0uyRqdImzPX2ADZzzBQnkyQIMX2crtlTXtKTZRaO5zWE1Sei6zl8qRSUltB2no
J1UvVLxRBm07SAV3p7Rf8F3zZ3ryuEt+QYmEwMAD+ZugpEQV2csD0NlV2HVDgSIuyjNDZZMezEOh
1Zuu4l4/2qMOa90hXGfg27fUqkgPcugvSy2d9rHC+RT/jFMrpcFLBjbZXJM4GxjvkEI5a1gHInIq
eiLAWl6aD1mvYmWU8LsfEtR8UoiT3J2UxMfxQ8EjElUbmjMNOa6vmK9c9u4i4sZ5qBUtPzcUY2Yp
/jrLk1Nh+fn+P/vVQY+IvL2P/mLqwWSIOOV5wWNLuVIptRNTHWPaYDEb2yHPsb5wFHbHRQiodA39
bxN63k91WpHu6crSNCxzF8SqcJJlHTtomwld3e1p1GVEtEy88OV953Ofp+Np4fymkXVWUKco+aPz
U3Gbi4enEZZBvpfyYLkyBBdSP15cMFyggQvKOFnsu4A8X1BxGs6Lo1xza3P8lxm1StdbO3Ecxly8
FbkDz0hIxNCLi7Lx9HPoDeDbjfkbMm+t0S/nAq6gVkJPnmeZtZPtlnouWSbTNTSh4y4MADi8Y5Gp
Jja/jaYH2v/3XeMpZs4HGfiJq7mnL2LAuuthMH1c+a48+fhRE7WVKt7js+3TOhJN2FoBO2cz/K2S
WND/+Q8pmqEP+PHvtScIJo5nyMMzysKAYwpundNjj1GVllbNMc5hyW8uvS/tVY2HkVl/NcLDKN6t
qDjgiFp7dDIEW33acM2z1IMKBOpZ0ikWWVi3mbMFRSabxgfWktuKWs6+kPDgXsmiVu+134XV6bte
F0DOodZsfQGzD5dgKe1/r6V/fxOgEYeCHd7YDI+yvkRhb4ao+XhrcKLqnsrRfjyhz51vCEdockve
dK2rz3GFOfKcpDRFj9BemM1ONpgTi4Mmo9wE3fZvSx5rI7Zk77eBvAw/ZUmpkcCmRImy9xVorzGW
Y9FLNZb8up5VI5ssxDdIFT7bLb27v8aNrhvuJieZcvMSnEAcZHWjUPJ7ifR8V+TrQkHc6R8uU20w
PVXnwfV3jXzQR8UbU+CS85bcd6S7Bl27AXQ75F7xJt/OU1qay2r47nyMP4jjAzEEoI46UtvAM1e8
AIcQH9uP0PUDNFeS/1FV1HWbp5HN7p9GWK2IbqU2t2QNz0rIIdKjxLulQtC02XF3OKXooQo51u5P
9nRUDI/Ut1ENVn+FTZjf+S09DkABz6uP1txLyV31Gv40FeSeC2hqzdJHAf9Au7pc5/78B9i8W0Tg
hm4hmUnyMUIxDIcgiu84dtdtvqtSCIyz4tPITSM0kZ3evrWQ6JbGmSWh5G3pRBXWV4D5HmlE3iWJ
pb/zmUWwn2J5oCn7zH4fFlXcLV9HFg73yI+sWTP8DOStDWD/pJzdnY7m1WHJAo5WlYHiG4qi2LAk
v1Q128jPvtiqxFMSS7EM3NqE5F3pT8sL3C7iUiCOwZpSKvfXrjsp3kK7MQRmrvRvc4OPUoaGXArf
9i3JD21TWpZuhXIx//RqH7Vi1eaDyH1myT52B/ZasVjQOP9+mowiNR2BF6cyEZ6mB9clLzBODNy7
5jS1eLCmNOQuBalc5v6NCt+gIAX6TvfSWP6O5GrGfyzNCKRseSu17uA6G0r9FybftDqHqNxxGBcL
Zg15JVtfSCYYpChSvDGBrh0F0lKHIKmWnwDQYWI3BTFKwEqH/HlSWXFTZ3L/yg0Fu0R2ShmTTGZG
4862z/qvkfTpfWLpQgvszNDORrYfjhCRRF0CQA3Jkb7bpP+eV2LaT1cHF0nNXdcBO5eiUYf6px+y
N6CIZKc9khlYGXZHxkPef5ZJ+fI+UPVIN6vE85IrRk7g+d00hcvIv5vMbfKbeedF2kyFXNF9BWPM
cm5N64YIunOwRFWY+zvc751O79838p5hmdQbBY5cTaiSeKO+uejAWZnaktCETWEd5vj8JLJK49ug
dWweb0tTrt/R5MLOacGNbzLL+bFn6w0gNjHly9kRXhRvvIp5j+W8Hy25KYRFaFeh6yxvl9LoiTyk
csMXOR6mE7eUkO3RTdqUHK0ZCpl0dizkjrKVM71OEg7dmY3twuRCcXZxuXbx94A05qpv5z7ZJrLB
gtB/SxleY6BQgWun2YqZzY10b6EykvKxl/oK8FH7ywSHNpKAVcEv/DLo42LSDj91OWMcUFObNm7t
gaG2B1+sKWLfMrvhdeFnRInlJJmeQRzShrRn7gDLrSM0zIqjQ/u87dxfz2Er/rN17t1xE2lXMnYt
IIZSkv4D5sv4q4B81MUoP95mNR0ZTPO6XRA7dP5d1sUmCUHfSHCihxDMG3ilZZqZuootZLvwi1qK
Iubjn1bDtD+WmsZXPU/XHgE3Bk+oMSeExwJObk+7kvZpHVNNDdUOoGyiSn3xFiGInZoBT3slxTFw
Uq0FzNfqlfcYZMjkM78iNaxeMOktxxk9hg86FdIcLr5M7byBEe7YlDlx0Z0aK0ODp1GALflvly1I
nF8Ka/L+6Ca6pGRBniX5IyL642s+E57XELrRTvP1YvuYLZBvenLIvKvEJErR6+timYG8lcW5YXcC
JUwtFc/2XZDaGb7smjz6CCvqmndeAFJDT71Ocp5SNvKd4qm9y2NjHqrrHsSAwZDZEsMMbkBY52WG
BVGnxgAGe1yeoXbBU/mc6o44qvn5f563OPzCeSC0LvTW9tyIrHcenVqxVB8bGHHJdN8kc1QBqnIF
b7O+s8NhWInt17JquKtcCfMFviyh+D0lHhuTRBtFWC+Vu0o17Xir0Hg5Xj6Dsp0Odl5i+OebFuj1
wG0GeSCEhJfOkNwEguQMtcLCFVmOIgvM7PFuzRzOBKNxpovS3JZ1HwI4+QKmdhKAiiRZc1zqpRSs
wTGaa7idV1kt2WxT9BSBCcQI6icreRqsTvKUCijS4UOmDXw/VEk0ltLG/KAqh3lKmEd1AP1924qc
1utO5jEiEFVxjNOo31UjJxdscIf3dQFKCSTMKyjZKyVtaaqtNqVGvnIVNIAdc6xaZGg1woHbt1yA
9O+tF9xW8C140IOywxyZqaKu/vcCgFn32qpd0lFbroc6lGKtynEZBqJTADel+TrkBa2lH9jvfJ1t
vei5Pt7qm3HI54ffSl92O237Id02+kjiozH562XlIPIYJZglA7LrywyrlG8nABmYDNgBD/7VmiMM
95NtDP7F0Y8Ip0Xp8I6p+3TfmKuToW+y7HmslmKGIELSPzJzSbKMdHAPKh7RQy8GSD3E4VWKFgrV
y0/GP+jH41KGRUS5jSeJgnZLWJ13xzXvN1sKUH8TXgC9CZhjcWWa5SNgpBFSTnI0BYYTpjuFZGJJ
LOXJ91YsH4ALM+eAT9u5AW4UXxaZBcAXuvY8SrpVcLIHuFSzFlbSNoNf7njXGJu5adOzPmG/eKQW
AaOakgw0NcmCj9sZIqnxAAG3yR+ZL/IAyfzpaxu09NmB+1GTjK2Urhski/RWHWNGX6aYV2ZBOmw3
SqGnnfo1Ffj7ubaUrisSILyv/WdZwyNLdvf8j5o9tJoxmN0bOvGzKB6wZ5/nqoNCyrEovbRLueX8
uaGMkwXbLjI8nC/GtGauoAVdP0QTNuTxEbKxBe7K4zLh0mdk3Jh1G2jewNpBG04VN550jxhkEw6u
FSZ9qlndDY4HZR21QEvvtNMbB5SWOu5JPGwfMi6wZMQezYE2gR+1XIQ46MZzrZeG2dDc/zDdKaEe
Qh/SBZ0boDV+mUEN17Jk7XVjs8dvgzLN5MHeVqkrYdtghBfeROeYQjVkah5bBYVJIu+7OEk0BQRW
6n+0sgn1Fu6agap3aTlo06r/EMO0qWauIZQ3at/KK/3zeBh00IhpWDznMlifhmRmwyLK8LsLTllc
xQMAiUVHRGnAfQvFYl10qVcwB1KXVaU2gi+hKeQZ5GlKKuccz5RnCf31b4BrCdzF7WPhkzNHKHAz
MJuTAMIVmoeN29ROkU3kdiRp/TcaoQFv+jJht8ysn/gj3CUNeQWYEWjPA+7Ur9XQLj/FuX+n3pq+
APBJ3DDH4sJMxDtNdRRsnVxX9cQScyD6oUEEPkdbK1V7PtEuRmd/1s5Xx7j1s3msCDKPd4Gale8s
18MMiWITC6wCq7sAf4SbndRGsPKDTVJOEBRZ0sZV5DzKsgG3elCfqbZhHNrckyM5YE9TJVEfI4vC
5tLjxQepme+2WhSq5oW1oXHB/862rXBqCR2b2FMox9OM16ykhw8y05V5iaiShXrGuRoevaQiz8Em
IhE7az1WWPPVb0MNji2uDkVjcQHGDDFcJPxj5nPAEJ2Q9oAPYwMIMg2XhpudyKW4GgiDkHZ/9JD2
Mmijxz/bZfmDSoPrIbRmNJtU55+phCMaUChA8CMYSaAjPoy8wMa7pezgwCzJMYoz+hfx8SjCqXfT
rooNJjTU+5selFVc0FjJKfDjqzaYi/3giLxks/Rc4CrN8QWQADBaU73JhbDFAgjnnH8Qbz8RWWxu
llBLdlp3Y7oP8Hv5S3lBrL/ek2BZYmmldIarNH/3cs+wWbO4OYtfE3pijqb7gQrRXujzYF6RASC2
Jdw3yQpL5IzOlixb+Vo+FfnYoVffn1EEfxApGhwBLeOznCGJujwZzSoFLsF6saOfl5ytOf1DSsnV
fBO4ZRRUvimBv6ZqhEbXo/H9OyNgWD7rep08rUeiISPedv8PHQGk7tX3v/7LpQCI/p7AUOZdCC4B
bzDAINfpAPVhs/1hX36dfd/SHzb3V6f3jS8NHgdp4BeXDtp+x8T0PQuanREPF01zDFBfXOwzK69l
L5yBharSOGSrO+R8umLSTxxxw4c3RULWvRcUFiJZplKuAJRGktuEv3W979Qot1Sa/s2+DKWzXqYe
poBZvvph6Xu7USPXOkQoVUaaNV3sstmlejOXlXtTqKHF9q1Wz7/PpSl/EOvE3J46zB3Fge5gvjqc
-- ==============================================================
-- RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
-- Version: 2020.1
-- Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
-- 
-- ===========================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity myproject is
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    layer1_input_V_ap_vld : IN STD_LOGIC;
    layer1_input_V : IN STD_LOGIC_VECTOR (879 downto 0);
    layer10_out_0_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_0_V_ap_vld : OUT STD_LOGIC;
    layer10_out_1_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_1_V_ap_vld : OUT STD_LOGIC;
    layer10_out_2_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_2_V_ap_vld : OUT STD_LOGIC;
    layer10_out_3_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_3_V_ap_vld : OUT STD_LOGIC;
    layer10_out_4_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_4_V_ap_vld : OUT STD_LOGIC;
    layer10_out_5_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_5_V_ap_vld : OUT STD_LOGIC;
    layer10_out_6_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_6_V_ap_vld : OUT STD_LOGIC;
    layer10_out_7_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_7_V_ap_vld : OUT STD_LOGIC;
    layer10_out_8_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_8_V_ap_vld : OUT STD_LOGIC;
    layer10_out_9_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_9_V_ap_vld : OUT STD_LOGIC;
    layer10_out_10_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_10_V_ap_vld : OUT STD_LOGIC;
    layer10_out_11_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_11_V_ap_vld : OUT STD_LOGIC;
    layer10_out_12_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_12_V_ap_vld : OUT STD_LOGIC;
    layer10_out_13_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_13_V_ap_vld : OUT STD_LOGIC;
    layer10_out_14_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_14_V_ap_vld : OUT STD_LOGIC;
    layer10_out_15_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_15_V_ap_vld : OUT STD_LOGIC;
    layer10_out_16_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_16_V_ap_vld : OUT STD_LOGIC;
    layer10_out_17_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_17_V_ap_vld : OUT STD_LOGIC;
    layer10_out_18_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_18_V_ap_vld : OUT STD_LOGIC;
    layer10_out_19_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_19_V_ap_vld : OUT STD_LOGIC;
    layer10_out_20_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_20_V_ap_vld : OUT STD_LOGIC;
    layer10_out_21_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_21_V_ap_vld : OUT STD_LOGIC;
    layer10_out_22_V : OUT STD_LOGIC_VECTOR (33 downto 0);
    layer10_out_22_V_ap_vld : OUT STD_LOGIC;
    const_size_in_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
    const_size_in_1_ap_vld : OUT STD_LOGIC;
    const_size_out_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
    const_size_out_1_ap_vld : OUT STD_LOGIC );
end;


architecture behav of myproject is 
    attribute CORE_GENERATION_INFO : STRING;
    attribute CORE_GENERATION_INFO of behav : architecture is
    "myproject,hls_ip_2020_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xcu250-figd2104-2L-e,HLS_INPUT_CLOCK=5.000000,HLS_INPUT_ARCH=pipeline,HLS_SYN_CLOCK=4.371125,HLS_SYN_LAT=8,HLS_SYN_TPT=1,HLS_SYN_MEM=13,HLS_SYN_DSP=23,HLS_SYN_FF=10590,HLS_SYN_LUT=132844,HLS_VERSION=2020_1}";
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';
    constant ap_ST_fsm_pp0_stage0 : STD_LOGIC_VECTOR (0 downto 0) := "1";
    constant ap_const_lv32_0 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000000";
    constant ap_const_boolean_1 : BOOLEAN := true;
    constant ap_const_boolean_0 : BOOLEAN := false;
    constant ap_const_lv880_lc_1 : STD_LOGIC_VECTOR (879 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_const_lv16_28 : STD_LOGIC_VECTOR (15 downto 0) := "0000000000101000";
    constant ap_const_lv16_17 : STD_LOGIC_VECTOR (15 downto 0) := "0000000000010111";

    signal ap_CS_fsm : STD_LOGIC_VECTOR (0 downto 0) := "1";
    attribute fsm_encoding : string;
    attribute fsm_encoding of ap_CS_fsm : signal is "none";
    signal ap_CS_fsm_pp0_stage0 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage0 : signal is "none";
    signal ap_enable_reg_pp0_iter0 : STD_LOGIC;
    signal ap_enable_reg_pp0_iter1 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter2 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter3 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter4 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter5 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter6 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter7 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter8 : STD_LOGIC := '0';
    signal ap_idle_pp0 : STD_LOGIC;
    signal layer1_input_V_ap_vld_in_sig : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8 : BOOLEAN;
    signal ap_block_pp0_stage0_11001 : BOOLEAN;
    signal layer1_input_V_preg : STD_LOGIC_VECTOR (879 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    signal layer1_input_V_in_sig : STD_LOGIC_VECTOR (879 downto 0);
    signal layer1_input_V_ap_vld_preg : STD_LOGIC := '0';
    signal layer1_input_V_blk_n : STD_LOGIC;
    signal ap_block_pp0_stage0 : BOOLEAN;
    signal layer4_out_0_V_reg_1620 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_1_V_reg_1625 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_2_V_reg_1630 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_3_V_reg_1635 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_4_V_reg_1640 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_5_V_reg_1645 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_6_V_reg_1650 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_7_V_reg_1655 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_8_V_reg_1660 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_9_V_reg_1665 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_10_V_reg_1670 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_11_V_reg_1675 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_12_V_reg_1680 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_13_V_reg_1685 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_14_V_reg_1690 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_15_V_reg_1695 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_16_V_reg_1700 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_17_V_reg_1705 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_18_V_reg_1710 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_19_V_reg_1715 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_20_V_reg_1720 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_21_V_reg_1725 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_22_V_reg_1730 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_23_V_reg_1735 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_24_V_reg_1740 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_25_V_reg_1745 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_26_V_reg_1750 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_27_V_reg_1755 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_28_V_reg_1760 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_29_V_reg_1765 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_30_V_reg_1770 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_31_V_reg_1775 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_32_V_reg_1780 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_33_V_reg_1785 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_34_V_reg_1790 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_35_V_reg_1795 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_36_V_reg_1800 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_37_V_reg_1805 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_38_V_reg_1810 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_39_V_reg_1815 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_40_V_reg_1820 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_41_V_reg_1825 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_42_V_reg_1830 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_43_V_reg_1835 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_44_V_reg_1840 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_45_V_reg_1845 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_46_V_reg_1850 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_47_V_reg_1855 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_48_V_reg_1860 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_49_V_reg_1865 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_50_V_reg_1870 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_51_V_reg_1875 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_52_V_reg_1880 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_53_V_reg_1885 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_54_V_reg_1890 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_55_V_reg_1895 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_56_V_reg_1900 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_57_V_reg_1905 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_58_V_reg_1910 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_59_V_reg_1915 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_60_V_reg_1920 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_61_V_reg_1925 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_62_V_reg_1930 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer4_out_63_V_reg_1935 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_0_V_reg_1940 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_1_V_reg_1945 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_2_V_reg_1950 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_3_V_reg_1955 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_4_V_reg_1960 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_5_V_reg_1965 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_6_V_reg_1970 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_7_V_reg_1975 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_8_V_reg_1980 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_9_V_reg_1985 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_10_V_reg_1990 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_11_V_reg_1995 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_12_V_reg_2000 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_13_V_reg_2005 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_14_V_reg_2010 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_15_V_reg_2015 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_16_V_reg_2020 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_17_V_reg_2025 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_18_V_reg_2030 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_19_V_reg_2035 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_20_V_reg_2040 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_21_V_reg_2045 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_22_V_reg_2050 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_23_V_reg_2055 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_24_V_reg_2060 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_25_V_reg_2065 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_26_V_reg_2070 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_27_V_reg_2075 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_28_V_reg_2080 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_29_V_reg_2085 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_30_V_reg_2090 : STD_LOGIC_VECTOR (6 downto 0);
    signal layer7_out_31_V_reg_2095 : STD_LOGIC_VECTOR (6 downto 0);
    signal ap_block_pp0_stage0_subdone : BOOLEAN;
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_32 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_33 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_34 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_35 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_36 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_37 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_38 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_39 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_40 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_41 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_42 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_43 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_44 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_45 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_46 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_47 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_48 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_49 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_50 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_51 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_52 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_53 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_54 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_55 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_56 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_57 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_58 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_59 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_60 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_61 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_62 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_63 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call33 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call33 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call33 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call33 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call33 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call33 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call33 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call33 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call33 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp11 : BOOLEAN;
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call163 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call163 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call163 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call163 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call163 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call163 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call163 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call163 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call163 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp142 : BOOLEAN;
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call229 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call229 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call229 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call229 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call229 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call229 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call229 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call229 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call229 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp209 : BOOLEAN;
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_ready : STD_LOGIC;
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_0 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_1 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_2 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_3 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_4 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_5 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_6 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_7 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_8 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_9 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_10 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_11 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_12 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_13 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_14 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_15 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_16 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_17 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_18 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_19 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_20 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_21 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_22 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_23 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_24 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_25 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_26 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_27 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_28 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_29 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_30 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_31 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_32 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_33 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_34 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_35 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_36 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_37 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_38 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_39 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_40 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_41 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_42 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_43 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_44 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_45 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_46 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_47 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_48 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_49 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_50 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_51 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_52 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_53 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_54 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_55 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_56 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_57 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_58 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_59 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_60 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_61 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_62 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_63 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_ready : STD_LOGIC;
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_0 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_1 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_2 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_3 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_4 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_5 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_6 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_7 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_8 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_9 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_10 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_11 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_12 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_13 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_14 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_15 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_16 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_17 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_18 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_19 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_20 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_21 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_22 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_23 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_24 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_25 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_26 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_27 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_28 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_29 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_30 : STD_LOGIC_VECTOR (6 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_31 : STD_LOGIC_VECTOR (6 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_done : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_idle : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_ready : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_ce : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_0 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_1 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_2 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_3 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_4 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_5 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_6 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_7 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_8 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_9 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_10 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_11 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_12 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_13 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_14 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_15 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_16 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_17 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_18 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_19 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_20 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_21 : STD_LOGIC_VECTOR (33 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_22 : STD_LOGIC_VECTOR (33 downto 0);
    signal ap_block_state1_pp0_stage0_iter0_ignore_call253 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call253 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call253 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call253 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call253 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call253 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call253 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call253 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call253 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp234 : BOOLEAN;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start_reg : STD_LOGIC := '0';
    signal ap_block_pp0_stage0_01001 : BOOLEAN;
    signal ap_NS_fsm : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_idle_pp0_0to7 : STD_LOGIC;
    signal ap_reset_idle_pp0 : STD_LOGIC;
    signal ap_enable_pp0 : STD_LOGIC;

    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2 IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_V_read : IN STD_LOGIC_VECTOR (879 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_32 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_33 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_34 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_35 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_36 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_37 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_38 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_39 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_40 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_41 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_42 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_43 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_44 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_45 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_46 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_47 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_48 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_49 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_50 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_51 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_52 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_53 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_54 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_55 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_56 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_57 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_58 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_59 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_60 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_61 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_62 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_63 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_32_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_33_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_34_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_35_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_36_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_37_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_38_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_39_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_40_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_41_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_42_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_43_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_44_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_45_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_46_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_47_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_48_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_49_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_50_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_51_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_52_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_53_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_54_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_55_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_56_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_57_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_58_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_59_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_60_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_61_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_62_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_63_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (6 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_32_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_33_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_34_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_35_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_36_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_37_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_38_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_39_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_40_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_41_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_42_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_43_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_44_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_45_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_46_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_47_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_48_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_49_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_50_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_51_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_52_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_53_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_54_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_55_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_56_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_57_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_58_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_59_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_60_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_61_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_62_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_63_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_32 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_33 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_34 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_35 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_36 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_37 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_38 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_39 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_40 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_41 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_42 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_43 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_44 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_45 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_46 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_47 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_48 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_49 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_50 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_51 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_52 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_53 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_54 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_55 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_56 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_57 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_58 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_59 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_60 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_61 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_62 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_63 : OUT STD_LOGIC_VECTOR (6 downto 0) );
    end component;


    component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (6 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (6 downto 0) );
    end component;


    component softmax_latency_ap_fixed_ap_fixed_softmax_config10_s IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        ap_start : IN STD_LOGIC;
        ap_done : OUT STD_LOGIC;
        ap_idle : OUT STD_LOGIC;
        ap_ready : OUT STD_LOGIC;
        ap_ce : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (33 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (33 downto 0) );
    end component;



begin
    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_V_read => layer1_input_V_in_sig,
        ap_return_0 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_0,
        ap_return_1 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_1,
        ap_return_2 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_2,
        ap_return_3 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_3,
        ap_return_4 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_4,
        ap_return_5 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_5,
        ap_return_6 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_6,
        ap_return_7 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_7,
        ap_return_8 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_8,
        ap_return_9 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_9,
        ap_return_10 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_10,
        ap_return_11 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_11,
        ap_return_12 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_12,
        ap_return_13 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_13,
        ap_return_14 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_14,
        ap_return_15 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_15,
        ap_return_16 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_16,
        ap_return_17 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_17,
        ap_return_18 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_18,
        ap_return_19 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_19,
        ap_return_20 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_20,
        ap_return_21 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_21,
        ap_return_22 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_22,
        ap_return_23 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_23,
        ap_return_24 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_24,
        ap_return_25 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_25,
        ap_return_26 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_26,
        ap_return_27 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_27,
        ap_return_28 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_28,
        ap_return_29 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_29,
        ap_return_30 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_30,
        ap_return_31 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_31,
        ap_return_32 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_32,
        ap_return_33 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_33,
        ap_return_34 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_34,
        ap_return_35 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_35,
        ap_return_36 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_36,
        ap_return_37 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_37,
        ap_return_38 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_38,
        ap_return_39 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_39,
        ap_return_40 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_40,
        ap_return_41 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_41,
        ap_return_42 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_42,
        ap_return_43 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_43,
        ap_return_44 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_44,
        ap_return_45 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_45,
        ap_return_46 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_46,
        ap_return_47 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_47,
        ap_return_48 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_48,
        ap_return_49 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_49,
        ap_return_50 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_50,
        ap_return_51 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_51,
        ap_return_52 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_52,
        ap_return_53 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_53,
        ap_return_54 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_54,
        ap_return_55 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_55,
        ap_return_56 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_56,
        ap_return_57 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_57,
        ap_return_58 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_58,
        ap_return_59 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_59,
        ap_return_60 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_60,
        ap_return_61 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_61,
        ap_return_62 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_62,
        ap_return_63 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_63,
        ap_ce => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_ce);

    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_0_V_read => layer4_out_0_V_reg_1620,
        data_1_V_read => layer4_out_1_V_reg_1625,
        data_2_V_read => layer4_out_2_V_reg_1630,
        data_3_V_read => layer4_out_3_V_reg_1635,
        data_4_V_read => layer4_out_4_V_reg_1640,
        data_5_V_read => layer4_out_5_V_reg_1645,
        data_6_V_read => layer4_out_6_V_reg_1650,
        data_7_V_read => layer4_out_7_V_reg_1655,
        data_8_V_read => layer4_out_8_V_reg_1660,
        data_9_V_read => layer4_out_9_V_reg_1665,
        data_10_V_read => layer4_out_10_V_reg_1670,
        data_11_V_read => layer4_out_11_V_reg_1675,
        data_12_V_read => layer4_out_12_V_reg_1680,
        data_13_V_read => layer4_out_13_V_reg_1685,
        data_14_V_read => layer4_out_14_V_reg_1690,
        data_15_V_read => layer4_out_15_V_reg_1695,
        data_16_V_read => layer4_out_16_V_reg_1700,
        data_17_V_read => layer4_out_17_V_reg_1705,
        data_18_V_read => layer4_out_18_V_reg_1710,
        data_19_V_read => layer4_out_19_V_reg_1715,
        data_20_V_read => layer4_out_20_V_reg_1720,
        data_21_V_read => layer4_out_21_V_reg_1725,
        data_22_V_read => layer4_out_22_V_reg_1730,
        data_23_V_read => layer4_out_23_V_reg_1735,
        data_24_V_read => layer4_out_24_V_reg_1740,
        data_25_V_read => layer4_out_25_V_reg_1745,
        data_26_V_read => layer4_out_26_V_reg_1750,
        data_27_V_read => layer4_out_27_V_reg_1755,
        data_28_V_read => layer4_out_28_V_reg_1760,
        data_29_V_read => layer4_out_29_V_reg_1765,
        data_30_V_read => layer4_out_30_V_reg_1770,
        data_31_V_read => layer4_out_31_V_reg_1775,
        data_32_V_read => layer4_out_32_V_reg_1780,
        data_33_V_read => layer4_out_33_V_reg_1785,
        data_34_V_read => layer4_out_34_V_reg_1790,
        data_35_V_read => layer4_out_35_V_reg_1795,
        data_36_V_read => layer4_out_36_V_reg_1800,
        data_37_V_read => layer4_out_37_V_reg_1805,
        data_38_V_read => layer4_out_38_V_reg_1810,
        data_39_V_read => layer4_out_39_V_reg_1815,
        data_40_V_read => layer4_out_40_V_reg_1820,
        data_41_V_read => layer4_out_41_V_reg_1825,
        data_42_V_read => layer4_out_42_V_reg_1830,
        data_43_V_read => layer4_out_43_V_reg_1835,
        data_44_V_read => layer4_out_44_V_reg_1840,
        data_45_V_read => layer4_out_45_V_reg_1845,
        data_46_V_read => layer4_out_46_V_reg_1850,
        data_47_V_read => layer4_out_47_V_reg_1855,
        data_48_V_read => layer4_out_48_V_reg_1860,
        data_49_V_read => layer4_out_49_V_reg_1865,
        data_50_V_read => layer4_out_50_V_reg_1870,
        data_51_V_read => layer4_out_51_V_reg_1875,
        data_52_V_read => layer4_out_52_V_reg_1880,
        data_53_V_read => layer4_out_53_V_reg_1885,
        data_54_V_read => layer4_out_54_V_reg_1890,
        data_55_V_read => layer4_out_55_V_reg_1895,
        data_56_V_read => layer4_out_56_V_reg_1900,
        data_57_V_read => layer4_out_57_V_reg_1905,
        data_58_V_read => layer4_out_58_V_reg_1910,
        data_59_V_read => layer4_out_59_V_reg_1915,
        data_60_V_read => layer4_out_60_V_reg_1920,
        data_61_V_read => layer4_out_61_V_reg_1925,
        data_62_V_read => layer4_out_62_V_reg_1930,
        data_63_V_read => layer4_out_63_V_reg_1935,
        ap_return_0 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_0,
        ap_return_1 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_1,
        ap_return_2 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_2,
        ap_return_3 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_3,
        ap_return_4 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_4,
        ap_return_5 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_5,
        ap_return_6 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_6,
        ap_return_7 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_7,
        ap_return_8 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_8,
        ap_return_9 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_9,
        ap_return_10 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_10,
        ap_return_11 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_11,
        ap_return_12 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_12,
        ap_return_13 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_13,
        ap_return_14 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_14,
        ap_return_15 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_15,
        ap_return_16 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_16,
        ap_return_17 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_17,
        ap_return_18 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_18,
        ap_return_19 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_19,
        ap_return_20 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_20,
        ap_return_21 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_21,
        ap_return_22 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_22,
        ap_return_23 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_23,
        ap_return_24 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_24,
        ap_return_25 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_25,
        ap_return_26 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_26,
        ap_return_27 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_27,
        ap_return_28 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_28,
        ap_return_29 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_29,
        ap_return_30 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_30,
        ap_return_31 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_31,
        ap_ce => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_ce);

    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_0_V_read => layer7_out_0_V_reg_1940,
        data_1_V_read => layer7_out_1_V_reg_1945,
        data_2_V_read => layer7_out_2_V_reg_1950,
        data_3_V_read => layer7_out_3_V_reg_1955,
        data_4_V_read => layer7_out_4_V_reg_1960,
        data_5_V_read => layer7_out_5_V_reg_1965,
        data_6_V_read => layer7_out_6_V_reg_1970,
        data_7_V_read => layer7_out_7_V_reg_1975,
        data_8_V_read => layer7_out_8_V_reg_1980,
        data_9_V_read => layer7_out_9_V_reg_1985,
        data_10_V_read => layer7_out_10_V_reg_1990,
        data_11_V_read => layer7_out_11_V_reg_1995,
        data_12_V_read => layer7_out_12_V_reg_2000,
        data_13_V_read => layer7_out_13_V_reg_2005,
        data_14_V_read => layer7_out_14_V_reg_2010,
        data_15_V_read => layer7_out_15_V_reg_2015,
        data_16_V_read => layer7_out_16_V_reg_2020,
        data_17_V_read => layer7_out_17_V_reg_2025,
        data_18_V_read => layer7_out_18_V_reg_2030,
        data_19_V_read => layer7_out_19_V_reg_2035,
        data_20_V_read => layer7_out_20_V_reg_2040,
        data_21_V_read => layer7_out_21_V_reg_2045,
        data_22_V_read => layer7_out_22_V_reg_2050,
        data_23_V_read => layer7_out_23_V_reg_2055,
        data_24_V_read => layer7_out_24_V_reg_2060,
        data_25_V_read => layer7_out_25_V_reg_2065,
        data_26_V_read => layer7_out_26_V_reg_2070,
        data_27_V_read => layer7_out_27_V_reg_2075,
        data_28_V_read => layer7_out_28_V_reg_2080,
        data_29_V_read => layer7_out_29_V_reg_2085,
        data_30_V_read => layer7_out_30_V_reg_2090,
        data_31_V_read => layer7_out_31_V_reg_2095,
        ap_return_0 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_0,
        ap_return_1 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_1,
        ap_return_2 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_2,
        ap_return_3 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_3,
        ap_return_4 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_4,
        ap_return_5 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_5,
        ap_return_6 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_6,
        ap_return_7 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_7,
        ap_return_8 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_8,
        ap_return_9 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_9,
        ap_return_10 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_10,
        ap_return_11 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_11,
        ap_return_12 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_12,
        ap_return_13 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_13,
        ap_return_14 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_14,
        ap_return_15 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_15,
        ap_return_16 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_16,
        ap_return_17 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_17,
        ap_return_18 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_18,
        ap_return_19 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_19,
        ap_return_20 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_20,
        ap_return_21 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_21,
        ap_return_22 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_22,
        ap_ce => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_ce);

    call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391 : component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s
    port map (
        ap_ready => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_ready,
        data_0_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_0,
        data_1_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_1,
        data_2_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_2,
        data_3_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_3,
        data_4_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_4,
        data_5_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_5,
        data_6_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_6,
        data_7_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_7,
        data_8_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_8,
        data_9_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_9,
        data_10_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_10,
        data_11_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_11,
        data_12_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_12,
        data_13_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_13,
        data_14_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_14,
        data_15_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_15,
        data_16_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_16,
        data_17_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_17,
        data_18_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_18,
        data_19_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_19,
        data_20_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_20,
        data_21_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_21,
        data_22_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_22,
        data_23_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_23,
        data_24_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_24,
        data_25_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_25,
        data_26_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_26,
        data_27_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_27,
        data_28_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_28,
        data_29_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_29,
        data_30_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_30,
        data_31_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_31,
        data_32_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_32,
        data_33_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_33,
        data_34_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_34,
        data_35_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_35,
        data_36_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_36,
        data_37_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_37,
        data_38_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_38,
        data_39_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_39,
        data_40_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_40,
        data_41_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_41,
        data_42_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_42,
        data_43_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_43,
        data_44_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_44,
        data_45_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_45,
        data_46_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_46,
        data_47_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_47,
        data_48_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_48,
        data_49_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_49,
        data_50_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_50,
        data_51_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_51,
        data_52_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_52,
        data_53_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_53,
        data_54_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_54,
        data_55_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_55,
        data_56_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_56,
        data_57_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_57,
        data_58_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_58,
        data_59_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_59,
        data_60_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_60,
        data_61_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_61,
        data_62_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_62,
        data_63_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_return_63,
        ap_return_0 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_0,
        ap_return_1 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_1,
        ap_return_2 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_2,
        ap_return_3 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_3,
        ap_return_4 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_4,
        ap_return_5 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_5,
        ap_return_6 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_6,
        ap_return_7 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_7,
        ap_return_8 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_8,
        ap_return_9 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_9,
        ap_return_10 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_10,
        ap_return_11 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_11,
        ap_return_12 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_12,
        ap_return_13 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_13,
        ap_return_14 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_14,
        ap_return_15 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_15,
        ap_return_16 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_16,
        ap_return_17 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_17,
        ap_return_18 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_18,
        ap_return_19 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_19,
        ap_return_20 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_20,
        ap_return_21 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_21,
        ap_return_22 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_22,
        ap_return_23 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_23,
        ap_return_24 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_24,
        ap_return_25 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_25,
        ap_return_26 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_26,
        ap_return_27 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_27,
        ap_return_28 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_28,
        ap_return_29 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_29,
        ap_return_30 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_30,
        ap_return_31 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_31,
        ap_return_32 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_32,
        ap_return_33 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_33,
        ap_return_34 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_34,
        ap_return_35 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_35,
        ap_return_36 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_36,
        ap_return_37 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_37,
        ap_return_38 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_38,
        ap_return_39 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_39,
        ap_return_40 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_40,
        ap_return_41 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_41,
        ap_return_42 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_42,
        ap_return_43 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_43,
        ap_return_44 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_44,
        ap_return_45 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_45,
        ap_return_46 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_46,
        ap_return_47 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_47,
        ap_return_48 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_48,
        ap_return_49 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_49,
        ap_return_50 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_50,
        ap_return_51 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_51,
        ap_return_52 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_52,
        ap_return_53 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_53,
        ap_return_54 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_54,
        ap_return_55 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_55,
        ap_return_56 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_56,
        ap_return_57 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_57,
        ap_return_58 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_58,
        ap_return_59 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_59,
        ap_return_60 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_60,
        ap_return_61 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_61,
        ap_return_62 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_62,
        ap_return_63 => call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_63);

    call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459 : component relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s
    port map (
        ap_ready => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_ready,
        data_0_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_0,
        data_1_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_1,
        data_2_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_2,
        data_3_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_3,
        data_4_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_4,
        data_5_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_5,
        data_6_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_6,
        data_7_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_7,
        data_8_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_8,
        data_9_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_9,
        data_10_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_10,
        data_11_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_11,
        data_12_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_12,
        data_13_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_13,
        data_14_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_14,
        data_15_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_15,
        data_16_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_16,
        data_17_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_17,
        data_18_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_18,
        data_19_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_19,
        data_20_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_20,
        data_21_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_21,
        data_22_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_22,
        data_23_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_23,
        data_24_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_24,
        data_25_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_25,
        data_26_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_26,
        data_27_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_27,
        data_28_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_28,
        data_29_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_29,
        data_30_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_30,
        data_31_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_return_31,
        ap_return_0 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_0,
        ap_return_1 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_1,
        ap_return_2 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_2,
        ap_return_3 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_3,
        ap_return_4 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_4,
        ap_return_5 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_5,
        ap_return_6 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_6,
        ap_return_7 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_7,
        ap_return_8 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_8,
        ap_return_9 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_9,
        ap_return_10 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_10,
        ap_return_11 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_11,
        ap_return_12 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_12,
        ap_return_13 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_13,
        ap_return_14 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_14,
        ap_return_15 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_15,
        ap_return_16 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_16,
        ap_return_17 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_17,
        ap_return_18 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_18,
        ap_return_19 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_19,
        ap_return_20 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_20,
        ap_return_21 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_21,
        ap_return_22 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_22,
        ap_return_23 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_23,
        ap_return_24 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_24,
        ap_return_25 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_25,
        ap_return_26 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_26,
        ap_return_27 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_27,
        ap_return_28 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_28,
        ap_return_29 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_29,
        ap_return_30 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_30,
        ap_return_31 => call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_31);

    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495 : component softmax_latency_ap_fixed_ap_fixed_softmax_config10_s
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        ap_start => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start,
        ap_done => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_done,
        ap_idle => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_idle,
        ap_ready => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_ready,
        ap_ce => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_ce,
        data_0_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_0,
        data_1_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_1,
        data_2_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_2,
        data_3_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_3,
        data_4_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_4,
        data_5_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_5,
        data_6_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_6,
        data_7_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_7,
        data_8_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_8,
        data_9_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_9,
        data_10_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_10,
        data_11_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_11,
        data_12_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_12,
        data_13_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_13,
        data_14_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_14,
        data_15_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_15,
        data_16_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_16,
        data_17_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_17,
        data_18_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_18,
        data_19_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_19,
        data_20_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_20,
        data_21_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_21,
        data_22_V_read => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_return_22,
        ap_return_0 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_0,
        ap_return_1 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_1,
        ap_return_2 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_2,
        ap_return_3 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_3,
        ap_return_4 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_4,
        ap_return_5 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_5,
        ap_return_6 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_6,
        ap_return_7 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_7,
        ap_return_8 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_8,
        ap_return_9 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_9,
        ap_return_10 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_10,
        ap_return_11 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_11,
        ap_return_12 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_12,
        ap_return_13 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_13,
        ap_return_14 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_14,
        ap_return_15 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_15,
        ap_return_16 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_16,
        ap_return_17 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_17,
        ap_return_18 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_18,
        ap_return_19 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_19,
        ap_return_20 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_20,
        ap_return_21 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_21,
        ap_return_22 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_22);





    ap_CS_fsm_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
            else
                ap_CS_fsm <= ap_NS_fsm;
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter1_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter1 <= ap_const_logic_0;
            else
                if (((ap_const_boolean_0 = ap_block_pp0_stage0_subdone) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
                    ap_enable_reg_pp0_iter1 <= ap_start;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter2_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter2 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter3_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter3 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter4_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter4 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter5_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter5 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter6_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter6 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter7_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter7 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter8_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter8 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
                end if; 
            end if;
        end if;
    end process;


    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start_reg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start_reg <= ap_const_logic_0;
            else
                if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter4 = ap_const_logic_1))) then 
                    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start_reg <= ap_const_logic_1;
                elsif ((grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_ready = ap_const_logic_1)) then 
                    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start_reg <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;


    layer1_input_V_ap_vld_preg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                layer1_input_V_ap_vld_preg <= ap_const_logic_0;
            else
                if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
                    layer1_input_V_ap_vld_preg <= ap_const_logic_0;
                elsif ((not(((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) and (layer1_input_V_ap_vld = ap_const_logic_1))) then 
                    layer1_input_V_ap_vld_preg <= layer1_input_V_ap_vld;
                end if; 
            end if;
        end if;
    end process;


    layer1_input_V_preg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                layer1_input_V_preg <= ap_const_lv880_lc_1;
            else
                if ((not(((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) and (layer1_input_V_ap_vld = ap_const_logic_1))) then 
                    layer1_input_V_preg <= layer1_input_V;
                end if; 
            end if;
        end if;
    end process;

    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then
                layer4_out_0_V_reg_1620 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_0;
                layer4_out_10_V_reg_1670 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_10;
                layer4_out_11_V_reg_1675 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_11;
                layer4_out_12_V_reg_1680 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_12;
                layer4_out_13_V_reg_1685 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_13;
                layer4_out_14_V_reg_1690 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_14;
                layer4_out_15_V_reg_1695 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_15;
                layer4_out_16_V_reg_1700 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_16;
                layer4_out_17_V_reg_1705 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_17;
                layer4_out_18_V_reg_1710 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_18;
                layer4_out_19_V_reg_1715 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_19;
                layer4_out_1_V_reg_1625 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_1;
                layer4_out_20_V_reg_1720 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_20;
                layer4_out_21_V_reg_1725 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_21;
                layer4_out_22_V_reg_1730 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_22;
                layer4_out_23_V_reg_1735 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_23;
                layer4_out_24_V_reg_1740 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_24;
                layer4_out_25_V_reg_1745 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_25;
                layer4_out_26_V_reg_1750 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_26;
                layer4_out_27_V_reg_1755 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_27;
                layer4_out_28_V_reg_1760 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_28;
                layer4_out_29_V_reg_1765 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_29;
                layer4_out_2_V_reg_1630 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_2;
                layer4_out_30_V_reg_1770 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_30;
                layer4_out_31_V_reg_1775 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_31;
                layer4_out_32_V_reg_1780 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_32;
                layer4_out_33_V_reg_1785 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_33;
                layer4_out_34_V_reg_1790 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_34;
                layer4_out_35_V_reg_1795 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_35;
                layer4_out_36_V_reg_1800 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_36;
                layer4_out_37_V_reg_1805 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_37;
                layer4_out_38_V_reg_1810 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_38;
                layer4_out_39_V_reg_1815 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_39;
                layer4_out_3_V_reg_1635 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_3;
                layer4_out_40_V_reg_1820 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_40;
                layer4_out_41_V_reg_1825 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_41;
                layer4_out_42_V_reg_1830 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_42;
                layer4_out_43_V_reg_1835 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_43;
                layer4_out_44_V_reg_1840 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_44;
                layer4_out_45_V_reg_1845 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_45;
                layer4_out_46_V_reg_1850 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_46;
                layer4_out_47_V_reg_1855 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_47;
                layer4_out_48_V_reg_1860 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_48;
                layer4_out_49_V_reg_1865 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_49;
                layer4_out_4_V_reg_1640 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_4;
                layer4_out_50_V_reg_1870 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_50;
                layer4_out_51_V_reg_1875 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_51;
                layer4_out_52_V_reg_1880 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_52;
                layer4_out_53_V_reg_1885 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_53;
                layer4_out_54_V_reg_1890 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_54;
                layer4_out_55_V_reg_1895 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_55;
                layer4_out_56_V_reg_1900 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_56;
                layer4_out_57_V_reg_1905 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_57;
                layer4_out_58_V_reg_1910 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_58;
                layer4_out_59_V_reg_1915 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_59;
                layer4_out_5_V_reg_1645 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_5;
                layer4_out_60_V_reg_1920 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_60;
                layer4_out_61_V_reg_1925 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_61;
                layer4_out_62_V_reg_1930 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_62;
                layer4_out_63_V_reg_1935 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_63;
                layer4_out_6_V_reg_1650 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_6;
                layer4_out_7_V_reg_1655 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_7;
                layer4_out_8_V_reg_1660 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_8;
                layer4_out_9_V_reg_1665 <= call_ret1_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config4_s_fu_391_ap_return_9;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_const_boolean_0 = ap_block_pp0_stage0_11001)) then
                layer7_out_0_V_reg_1940 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_0;
                layer7_out_10_V_reg_1990 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_10;
                layer7_out_11_V_reg_1995 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_11;
                layer7_out_12_V_reg_2000 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_12;
                layer7_out_13_V_reg_2005 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_13;
                layer7_out_14_V_reg_2010 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_14;
                layer7_out_15_V_reg_2015 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_15;
                layer7_out_16_V_reg_2020 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_16;
                layer7_out_17_V_reg_2025 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_17;
                layer7_out_18_V_reg_2030 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_18;
                layer7_out_19_V_reg_2035 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_19;
                layer7_out_1_V_reg_1945 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_1;
                layer7_out_20_V_reg_2040 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_20;
                layer7_out_21_V_reg_2045 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_21;
                layer7_out_22_V_reg_2050 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_22;
                layer7_out_23_V_reg_2055 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_23;
                layer7_out_24_V_reg_2060 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_24;
                layer7_out_25_V_reg_2065 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_25;
                layer7_out_26_V_reg_2070 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_26;
                layer7_out_27_V_reg_2075 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_27;
                layer7_out_28_V_reg_2080 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_28;
                layer7_out_29_V_reg_2085 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_29;
                layer7_out_2_V_reg_1950 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_2;
                layer7_out_30_V_reg_2090 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_30;
                layer7_out_31_V_reg_2095 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_31;
                layer7_out_3_V_reg_1955 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_3;
                layer7_out_4_V_reg_1960 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_4;
                layer7_out_5_V_reg_1965 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_5;
                layer7_out_6_V_reg_1970 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_6;
                layer7_out_7_V_reg_1975 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_7;
                layer7_out_8_V_reg_1980 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_8;
                layer7_out_9_V_reg_1985 <= call_ret3_relu_ap_fixed_ap_fixed_7_1_0_0_0_relu_config7_s_fu_459_ap_return_9;
            end if;
        end if;
    end process;

    ap_NS_fsm_assign_proc : process (ap_CS_fsm, ap_block_pp0_stage0_subdone, ap_reset_idle_pp0)
    begin
        case ap_CS_fsm is
            when ap_ST_fsm_pp0_stage0 => 
                ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
            when others =>  
                ap_NS_fsm <= "X";
        end case;
    end process;
    ap_CS_fsm_pp0_stage0 <= ap_CS_fsm(0);
        ap_block_pp0_stage0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage0_01001_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_01001 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp11_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp11 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp142_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp142 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp209_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp209 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp234_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp234 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_subdone_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_subdone <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_state1_pp0_stage0_iter0_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0 <= ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call163_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call163 <= ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call229_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call229 <= ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call253_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call253 <= ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call33_assign_proc : process(ap_start, layer1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call33 <= ((ap_start = ap_const_logic_0) or (layer1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;

        ap_block_state2_pp0_stage0_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call163 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call229 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call253 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call33 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call163 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call229 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call253 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call33 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call163 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call229 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call253 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call33 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call163 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call229 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call253 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call33 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call163 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call229 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call253 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call33 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call163 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call229 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call253 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call33 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call163 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call229 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call253 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call33 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call163 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call229 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call253 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call33 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_done_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            ap_done <= ap_const_logic_1;
        else 
            ap_done <= ap_const_logic_0;
        end if; 
    end process;

    ap_enable_pp0 <= (ap_idle_pp0 xor ap_const_logic_1);
    ap_enable_reg_pp0_iter0 <= ap_start;

    ap_idle_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, ap_idle_pp0)
    begin
        if (((ap_start = ap_const_logic_0) and (ap_idle_pp0 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            ap_idle <= ap_const_logic_1;
        else 
            ap_idle <= ap_const_logic_0;
        end if; 
    end process;


    ap_idle_pp0_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_enable_reg_pp0_iter2, ap_enable_reg_pp0_iter3, ap_enable_reg_pp0_iter4, ap_enable_reg_pp0_iter5, ap_enable_reg_pp0_iter6, ap_enable_reg_pp0_iter7, ap_enable_reg_pp0_iter8)
    begin
        if (((ap_enable_reg_pp0_iter8 = ap_const_logic_0) and (ap_enable_reg_pp0_iter7 = ap_const_logic_0) and (ap_enable_reg_pp0_iter6 = ap_const_logic_0) and (ap_enable_reg_pp0_iter5 = ap_const_logic_0) and (ap_enable_reg_pp0_iter4 = ap_const_logic_0) and (ap_enable_reg_pp0_iter3 = ap_const_logic_0) and (ap_enable_reg_pp0_iter2 = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0))) then 
            ap_idle_pp0 <= ap_const_logic_1;
        else 
            ap_idle_pp0 <= ap_const_logic_0;
        end if; 
    end process;


    ap_idle_pp0_0to7_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_enable_reg_pp0_iter2, ap_enable_reg_pp0_iter3, ap_enable_reg_pp0_iter4, ap_enable_reg_pp0_iter5, ap_enable_reg_pp0_iter6, ap_enable_reg_pp0_iter7)
    begin
        if (((ap_enable_reg_pp0_iter7 = ap_const_logic_0) and (ap_enable_reg_pp0_iter6 = ap_const_logic_0) and (ap_enable_reg_pp0_iter5 = ap_const_logic_0) and (ap_enable_reg_pp0_iter4 = ap_const_logic_0) and (ap_enable_reg_pp0_iter3 = ap_const_logic_0) and (ap_enable_reg_pp0_iter2 = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0))) then 
            ap_idle_pp0_0to7 <= ap_const_logic_1;
        else 
            ap_idle_pp0_0to7 <= ap_const_logic_0;
        end if; 
    end process;


    ap_ready_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            ap_ready <= ap_const_logic_1;
        else 
            ap_ready <= ap_const_logic_0;
        end if; 
    end process;


    ap_reset_idle_pp0_assign_proc : process(ap_start, ap_idle_pp0_0to7)
    begin
        if (((ap_start = ap_const_logic_0) and (ap_idle_pp0_0to7 = ap_const_logic_1))) then 
            ap_reset_idle_pp0 <= ap_const_logic_1;
        else 
            ap_reset_idle_pp0 <= ap_const_logic_0;
        end if; 
    end process;

    const_size_in_1 <= ap_const_lv16_28;

    const_size_in_1_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            const_size_in_1_ap_vld <= ap_const_logic_1;
        else 
            const_size_in_1_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    const_size_out_1 <= ap_const_lv16_17;

    const_size_out_1_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            const_size_out_1_ap_vld <= ap_const_logic_1;
        else 
            const_size_out_1_ap_vld <= ap_const_logic_0;
        end if; 
    end process;


    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp142)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp142) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_287_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp11)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp11) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_281_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp209)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp209) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_355_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp234)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp234) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_ce <= ap_const_logic_1;
        else 
            grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_ce <= ap_const_logic_0;
        end if; 
    end process;

    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_start_reg;
    layer10_out_0_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_0;

    layer10_out_0_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_0_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_0_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_10_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_10;

    layer10_out_10_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_10_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_10_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_11_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_11;

    layer10_out_11_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_11_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_11_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_12_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_12;

    layer10_out_12_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_12_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_12_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_13_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_13;

    layer10_out_13_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_13_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_13_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_14_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_14;

    layer10_out_14_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_14_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_14_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_15_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_15;

    layer10_out_15_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_15_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_15_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_16_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_16;

    layer10_out_16_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_16_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_16_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_17_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_17;

    layer10_out_17_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_17_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_17_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_18_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_18;

    layer10_out_18_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_18_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_18_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_19_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_19;

    layer10_out_19_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_19_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_19_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_1_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_1;

    layer10_out_1_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_1_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_1_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_20_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_20;

    layer10_out_20_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_20_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_20_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_21_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_21;

    layer10_out_21_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_21_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_21_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_22_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_22;

    layer10_out_22_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_22_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_22_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_2_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_2;

    layer10_out_2_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_2_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_2_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_3_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_3;

    layer10_out_3_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_3_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_3_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_4_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_4;

    layer10_out_4_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_4_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_4_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_5_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_5;

    layer10_out_5_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_5_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_5_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_6_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_6;

    layer10_out_6_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_6_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_6_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_7_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_7;

    layer10_out_7_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_7_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_7_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_8_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_8;

    layer10_out_8_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_8_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_8_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer10_out_9_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config10_s_fu_495_ap_return_9;

    layer10_out_9_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter8, ap_block_pp0_stage0_11001)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001) and (ap_enable_reg_pp0_iter8 = ap_const_logic_1))) then 
            layer10_out_9_V_ap_vld <= ap_const_logic_1;
        else 
            layer10_out_9_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;


    layer1_input_V_ap_vld_in_sig_assign_proc : process(layer1_input_V_ap_vld, layer1_input_V_ap_vld_preg)
    begin
        if ((layer1_input_V_ap_vld = ap_const_logic_1)) then 
            layer1_input_V_ap_vld_in_sig <= layer1_input_V_ap_vld;
        else 
            layer1_input_V_ap_vld_in_sig <= layer1_input_V_ap_vld_preg;
        end if; 
    end process;


    layer1_input_V_blk_n_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, layer1_input_V_ap_vld, ap_block_pp0_stage0)
    begin
        if (((ap_start = ap_const_logic_1) and (ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0))) then 
            layer1_input_V_blk_n <= layer1_input_V_ap_vld;
        else 
            layer1_input_V_blk_n <= ap_const_logic_1;
        end if; 
    end process;


    layer1_input_V_in_sig_assign_proc : process(layer1_input_V_ap_vld, layer1_input_V, layer1_input_V_preg)
    begin
        if ((layer1_input_V_ap_vld = ap_const_logic_1)) then 
            layer1_input_V_in_sig <= layer1_input_V;
        else 
            layer1_input_V_in_sig <= layer1_input_V_preg;
        end if; 
    end process;

end behav;
c5+KFGFaw6XTh5lgXq+mnhUtX0Tx1xNvHmttdB224JT71sTXO+zB9OtReqfd4I0Foh+DnEamPd2c
kP2KrpMMo1GlGda0BH2IHbj1COH2yIGKmjZPqNSgmTbvpKhc68IOCUcOkijBFek3OWCM0b5wZHf0
CfNNMb/TtGyriYGKNjHDNVQUWmmerae9iNwWZz1Ed3hEuL9DrIhhU7aPLEyL9jxqrcuw1zxqCMAy
YTMdlnfcj+10lTFwovNreBFE8IoJbpo8dYN50FgUgAH8PIRq/w5PHvxluW+PiSZYuraOXzurvlGn
61SWuPmvDSIZzIadRCS7We2wl9gz9uV+SkFlikDHhljZ2LcWFdbsSAf2jvRiaBn2c+MyaKbbEQG1
vjJcRumhZalWIDT0tF/E0KWaaO1+4cxCi/7068BJ+lu6IilyHJwgZtjU8yBfXEoSb3OsCUT9LhQG
rNBn1M1ajN+EoTzG0+4CfS0sFys1dOE50r7RZ1YdsoDozBoVkNAcoRuLiAEHeyAFASGKJ3EetpSV
ezMdmESglxo5gCJ9+0BxxmYzkCQr7zWZxR4osDSFA4JtW2riUDV5sCxmfI+Fr/SmnLYE5u/3U3es
ww5RxN/XckgjMd3voHcGgGX7VcKw0D+lh4Gs5m+s+B8dDZkI02vZg54mxOoZbxyoktH2TX6EOHv8
TZQv4wB50dF3EZqxV6yUz/JckvNo8xw0cJZI29z3yYinQpRtZHS/OOAO3lxnLcAbjnaasN0EFI2/
Bjzk6U/RLl1j4EicRrZ7MoUKig6T5JViUTw+I8JRWF3yF2NMdDRLNSRJbbYPn3AaBXV5xFg2kAbg
ZzMWsAMkLojLIC3N86bb/4jNKWV1/IUz1ggbY3D17XPUX6m9/DGhCmdIw3Gq5IzAp1kHwAai4ZI7
dm4rCBG2LFyNcfyKMyodMCBiJ4jTvItwvcb7eNhaFuvaqjtf3SVVtxvHZOpFUAzrhK+U4C2rsDmM
6ejdoOiqiaNGr5iedrD0EhSq+7NOCjoXy6by9jDLe09eGzcJiXe+4QE8WWYFvePrvCtqnJ/a1CeB
NPE3/NwisgSYDOesZgPeFA3bpiwcUDIQ0LS4kvJ2mQdJRaOEZz0sILP1bvRA87iWKRPrUMz239yF
ANpFM3LGU8gpcGBP2iq8lhIWm2sfqC++ZKWGVLdM/yAAgfY33vaEHDK+c1y07tkibidiod9iYKWw
gbKrJaKFlndYH5v4KmXn5j32AD29yh0nvgQYPebJmBrsb6cbrktu8tCeOeVT84LVb57FykNHMrwq
4+xEjhttXfaZTK8tiMVmFLiTy+TAtWie2PTXxmRDcS0kBeQnTFen3Hudr7HRsJrT4mcwqxJKT1oy
Pa6sGKJpBJfUAFLE0mRZ/2ApA4XT/YzUBxFDkpk40dl6bPDpyy6Z6vWE76/noMpNgB/mlQg1jG42
g0KhjBJhDq0kT1n/tpf2yLGT85USilw6/8M0s6urB5+ThQy/SGrrnt5Q38m+hVhSYMDSJ6pqb6RC
OxhvoMj4sUTRN/W10BJ63ErN+a4UmvIT4xRMFHKpyNW06cVvhBgOrtymHb32CeFjDZRZ2NDdBAsQ
AvT5bog0WQhFIeDJle0iQ2QZ3Rtmc9/0BnV72QGiets/xokTxyVoLLbavE/W72t5lEd0salF1TzF
weUyLhursgLw/z57cTac/FS5SGKfFQdm3RzTusn8Tsxs7eqsvikIaEL7u87gQ9PBF+llLNWFl94K
VL5LN/p0kSgg+YL6DAms+JqSVXjaCbjRjM0brn1z0kUMKyzaTB7jNOf3m8uUKAExnfnyc3h0uQxM
5hefRBb00kcc7KC0Sa8aDQ14vbO0mCeZRQXELFDA1ANiOtt2dHvqc7OUaS1c7rPyt9AkIlaWn/St
YDMs6qm5YXw5XULvweSn+vXx+5MNBv/CPhvxpUJbY76emuEhuhedYD8+WzH+I9sS85voiblqmzOu
RKH2RCHUcTqdj7AlOR6CAkUvK2RmH3uqp7JhTAuxw69RUj4GyBLmoVOkD/z6MYB7dyyBGbSrhdAY
SyF1oqjG8lFcMNh5ESM1cMuh/eXmsUJ43o0Lqfc4j8UnNS6z6vjUTNUcPbQdiVf9gwGCr6l6fUQx
1URyke4+Dtud/W9NQWkDCL6wgTURH2iDvvcciG4R0hjXIIO7KJC1NA7zWJl5TR1rdND2RoZfzJue
A1YWYIxLOhTKZdXdhZqxR2+c6SLmqTxsiZO214106/OZ5KNaiBtN+KFFP8k0HxITYOMtw2cE+woc
guIKBKWHyStd7KpxKsDGboZOR1YoUHg7jWiTvEVG+d0DIp5CPQnv+mZq4In/pVu8voqi5MYcyinT
YLsk9UsYBVMszPA3RWbQEAUpZP9NL0zprKiCTaHJg2Xwm/zay8GxKP++La44FMwuNCNlwuLndNVY
l+uMoq2LWvThXtt3Asf8Xf6KWYyt6NPlAd4BgQzsJLVLmSOwJSBVlPd5oGA5f5cpIMvxeZw1O3fh
hDQ5XkiYdCHVlB8sLS1uovtnLw+muJNpBabC+Fyw9IbQ0xRc17On2ZRDjvwuIWE13RJPksGTcNuH
WY1CvbZYo1Ace4blOVoO+p3IbcTbInxjLLIJoZQURuPMSRAy31pfODxor6wBP3Nlk1l1sxBSF5CR
PCdBbeVh8BGG/bL4J3rEobRRgmVhinycNnyKCEal5I1avS8s4SaA3cvSSS7rHBZFvv7PChuFbYF0
h20vDzSFy3598z//u7MF4ZtQKmKB8WoIokWwMYc2hRnXEIWlgHNy8kU43npqHuPXrhKWbiMIVFBT
5o8ZcQZBoa2tUsbur29x4/VS4dYQ7QeuiSwKIswaypZT/JlEJrWi6smbCjbAK/4Og9rSEp7JqvA9
vKWhA/cAsu1gcBArx2uwaUQe07tcMMJB6hIvqbBF5UFAz7qLvgBQhhv/LF3xD1CoxYuqh9km0GwW
pvrrE9fwVCw6Jk2UjpCy+h32UfhozAwe87fgoGGsIR2y798KKhmjcDCcOakc5oW/noWAYOJ8OamZ
kVNICUdygvtPfQP2vn1kmn+H1SUEBfXAC7OeU5N7mozMFx0ckO8UuFWrTSQ7XMt+axSlBaq8oL5q
P2mWbVvPs1f28UUU3TraJDneVxp6YzVVC4jnQ6Gop0CJcNhaU+iMaJxiCOiwFHJcRL0SDdTWDFJ8
NDjFrwlImbHgnnCnImylUWHqHdg9r3LIThUordUj4v0zM2iwcKttRxdcMbr5AEoZjJCwjtj/ewhU
eLvjGH6arBMYuC7aZ0l2O8tu46KrQCiNVRg50TqzYVSsQ+0EYGre3L7s8KE1eX6o9YhSYO8hi1b9
k0bLssRgpCkSaVqX1Kb86EzeTCi3hSM+JAQXnba7M5q2vP69Hv4lbXDCPO2nYVGTmNYQham3iAXi
SOL609gCiiVCK84hejMgVoqPD3aEfxwmpFj2O4Kea4OCwn+/TZmqawSmDYSohaL++uYxcGEbYRda
pn9S89KCQztuwCvtP9v0/rBjMxcG7bkUvRezE+i8tvDB4/4fPGLFEcVDfs8BLTMKZyhmA29GAzIq
kL0ZAWQYCuSFo8VHgt/DPbKMS4LbZwshiI/clq9HylcTEY5XMDLG0LAaYSju3lW6Wi/DIc/nZAr1
u92u8Ap3kaBCgf+vhcn3NBxHe3bZjKB2879dAkP1kbFd/5RSNLTc+/Mu7Ab7v+atToWQY4E60ljY
P6AD/Xut7Ettb3DNGdp+DyJNjMjo2EgWjIOi882GEO8WRMO1MhHFyu9uzxZ+107cHeSFTAKcqZRB
dH/wXVxexMnHfNlnqbaZWp7/VW7CTy0Z6msxfNbi1QuzYJjOXeY4DB+WRT4AsJQUaHxQAPcXmRoy
ZDV/uIo74zFzlTJ4t9m3HQboLg2S+LMpSmWnudQ4dQJnb/dufs12Q9C22A0TIXyybkas2f9mQYPz
IwWNjcnmPLiTPdC6Xg39XX8aIcaNPXoKKggWTKe4oliytoshNHBQsv6tb8fjhMDsxJQOneqJq6Hg
Vlk8Fhv44u91llIljo8Ni7O+3YHGljeCj7BeilojmcBJyoW5A/EZ4xqEsT/iAZIik9jPckxdAjSu
rZiS5EIhlIKGFp4DkW1ASKjED/kYaNaaJxVYo7ePeg3Cq7/2Z34Sm0fMfra9HqguxfocwadW3X5Q
eP2MKyLUwP+sDXp8uWzLmh0JRHOAtN7VKn2F95A2cYdPnjSYGGs4C1vAHHt8vPcwb8UNrH5dfpYK
Au+4UJQAK8rUHDAIdxIRhVOFHnmDEOwd0LA+zxNwh+HHXYtbkKMXCZtr8+C1cvtfGsZhtn457zPw
W5q2d58Sg1j5Hu1fPZox3Qq8d7OCKPUXeCreJFrXhgYmQiNktwc7vN8OWnMNV/ywP9ocNI/ykMfV
rCLK3FqVQGZm5tY3xsgPDsi3OlrlYRoQZPMdv2feeWf4znaH4XJx0o3tndd35VDUJ8qup7IAABFR
1OaEoMrDd8uDfIVJszTK7z2i2M2OIk9pr+wgzXY/r4uoF7qfOW9x/F9beTudzWv0qC8Gi0qQh6If
BHtkULcMQH81QEBIA2DLytyPeS5qmkI/xQAG31kcytTPu7l9slNf5q7BZmBKamn0BuB5/1XmwR9l
tjp9Ixmi1b1XOcqdwDf7yIVzu+oeEYRBUamo0M7R10XKxXIaRxeKeUwMOBTvumNsMbMbc04BOb17
Lx8P1o2CPLhj6aiJ0kQJAPtmZ9nrXQl7PBiZS30Nu2imt4DnL4CNQTcc2jMR0haYvTRc9r86RrRJ
YUWiDEJj9yGX838GMYun3qxzx92TtXdJpTuSR3oFzfrqMVB7GUrR5KF/685cVcJzsxGCghEPl64a
Xy70ZNKYrD8vWaHDhvylLAy3OjN2quu9l5PW7VU2FrBAWw1eWQjZb20UZRLghc3pjpz1pnAfJHxR
Kx9/H9KSP/0CiP3g1kQag+DMQ9u7odhbYoffYgC6d00IucatqUpzKCwYd1CCIu2lEd+/DG9rBdqm
Xk7DpMf8bXqIym8Hy4OzT0xXkqs76xKS+f7XPW0iKxFcFFnL4PtYJnONQd1CJX0eUjroJ6GVzY7Y
39quLdKJo7FqSzdLGCTlMZwr3y39N8vqsRQeVqkxI+cQMol0CG3ttAojuaVzwn6B1lRm/DQyDBhy
SUDpgbD50+klsUTDZcq+ZscMpZaUkTt3xYsnFjwv65J/EQ1YorNUF6N8joVIPYNkKyvFGovSLlIn
3bNEbGi7NWe7U2z6wUqQI0Xy/RG2BLhigYUGn/su0mEKLx93lBMEcBAoFfZ5r1FcNeIndrHOXYGA
Ofj5BIQef+RycG/Iec3CatPSKuRz4q5ciC7HTt9H0IAREcHiC0qyw/abe4QarXvqLkb9uvdbihGt
U3BiMcKoVBsQWHtxeqvbo2wiD15Xc1gJCUjA3KsOB71QSEjeC6buVVvioTT8NEAA4FZ7CkQ87qgs
2QlqlWe2YuW6aXagGLqgj2lPBAK+b9HYt+iGlJzrbLRj0OAYQU3kGlvKTCvXxymZxrlGA28/bPci
uRnVK/ofVDlyU4g9+gn4YrKGUKN/Swx2UGI+FPrMkSRGwZKQLpmTb9UOv59uCuDwh4RYVRytu6LR
fpjysSOX47uu1fW2srC5XIhXOCP5GynlXqr41EigMV2CZ5fFtxh9rij119l8IcYm62Agyl9Cs86E
1uEiBHox7iOpHcDVkeqmFT3DrsUhOoWKsshmoOpm1GrTe4I5iF/t+sdhiXRxZoDtk1dU6++ObN03
+GVdrsyGGxu07PrEWzHFxyMZ9+l/B8Fp9u1HH7kfjqt0cHpI+l7MzM9Ehu4ErG7vSgf8F+hLLEVU
P2/Pm1WOCpeNCygSIFS7Ts0Y+tCyRvfVziAIgdDETSCVcjeF3JTeR24dzWr5OVqOSxuvfnxsAXml
TGy/6jSHkNijSrlc1KSJcrVbtifKC0n07hmVrVWkOoQin7lIwbvr1S3FmBM1W16jtbKU5Z0RH7dW
i7k0N0onpw3+sYzkyEx8ozzsGSHIFB7uDbBfxG+LJz1/NyEA5k34SYt9R53bPJjThFsCrG54Od6x
3mxbajHj2BlTk+mDHCC3aDwTVu11zjsr5Eg+zd1XbBYlcgIS7UO9hOUdYGmdOP8qWq9DUI+Qtn9i
xLNbAPwLbnPbTcnCDWgGnHF2TTkLatFPFsaw3nCYA60tyMioy10He6xnKIIH8YEc9bLE5nSlWwfg
Iwr5NB3NsBiRx72D54du9h+usjApsvCAbURhS5ScPCm0F/ioS2YQ/r5KrotL4s0IsMnl1JNunOR3
ypXqMVtKxfqLtDMATW0wSo6yrNLlzkaIDUsub7hYJh74vymrLMBCZ0sAqtOWhQHF5AWdiN3Ju0nE
auJx80XSQnZrf3txup7bONYLtrIf9oO2KTRrPx8acGX/QXCpM0gR0KUKg/DREf8NrVdvJXV814pA
OFGA7UM3omtllacGqom9pDohApobQIHHgQ0Vm8ClJWW6U18Jw9MBrm02zXjrd3Zolds8k7GAIcDS
vXyNcsp5Fj84hHn/lK4VdRqM51hl9UMVRT7DN0CQJktjrpYEmEtbUMqcYx0jRRytwzCAz9n4LZzz
MYHr5mrYmIhJjmB4M7onELdC7fDwBsEzW27poGMMmwy8TYA2bM0LQT6xUmb/ohwJ+TE6/CEaLYZh
rJlsjO6YvkelV89f9PGJPWu2xBaE3ohMv56aBdSYxKqpLgaCHINVTr7/m5FFcU2R5x9vG6ZrWtKH
IlXltquxTHDuD6bliu7qsmayM13V9U93N4mJoT3qhUjI1/r5ZRDd+QaV+Tr4lJdGCagGdJ+xJWXM
+wJbQJiOAQws8TFgNYAae2+kh+3sFQVwj+n7NA+c3vnzH+sQclrwlu1OzaMGwNZetuuc1CfWWM0i
hVSsvzNWc6aEyra9MJO5aVdkKna8Ymi1nzJjHVrVok54JFGctBdQbPij1wVePqH5cqO0zCQy4Ey3
hbTYDNpjzy3OrVO67rPxVMouwlmznKJTmsqaL3bMbUG+GfBeNKc5DxophzIUE4D0ZTMx7KtRvoFa
lfzBI18XMLeZK5FOkVtcT9GL6oAeqPcrpOBdivTWBgW/M2mNeNw2PToZ82WXyK1m9TFoH2i8ZOrW
m6xiZ3LxWc0IBC7HPCAkYD0oBs/+aRkyi4otCE8ouYU/sh2CPg7ur4sDRyrbYgLa/3dn/prwmIQi
X8xiJOiV/Vsmfm9foZbObS25D78FsrNLXDHnfiZ+K591IkbLO6xntLpd/4F0GoqOCwbPgnncgUPd
R47NBzbVwEOz6hunI3yla069NU9tkpcDbXXmpNNpunjLrMGdmpq3cXr7zMOZdbCJH558tvsYvdOj
992acpIT/vRa0Qk/AXpi47LBm9VLnqfT5MfTsQN3sHwca9mP3ZsgyUTdRsGKuCveZkPAJeDui05e
YN8BYA7sxuRUVxQ+gJ6UaEeRI6TJx2yYguXbD3FRid5YcNnyPdhmfa4gsE+35G7EpINg3WYG6LDn
RscT4YHFVJ12CWWy+yGVJoOWx4qA6yZTwCWk4roqlmlq7yGeyssrRHqDGcwtO7P+7H3RUqInMYT8
m8OygsZIbI6ZgkT53/f8YQ2oNsKmV95wORHAr4XJyxyDNTYQjPZYwT6liYMw5zrn7lN+YBZR061Y
AsL/Y6jk0Rs9zuv8Kvfdf/g60n6PRhlFb4XBIwc5UlBYfgzZrNhkBVmwtBjcgABA+GI/tHPbeCK6
/aIxRIJLNC2xfHQ22pSjrv18gqqEM0bNbJXIYya98ogu+LnrK7wPSQO2IqqVElryLkAtF9Z/CX/o
ADe1WqJnZRPqDAE5ugHCmxoM1EJuiASbDxqAQYC0WJC74iKFp2NXYFNdT5dclKv180NS3YV4LVGS
LeB+dbMPMy03ud7UnxYLW/VcP5unG20NQsUm8J9nEx415Ox/asEDZRL319D4Tpv85Aoz+Vd0bWI/
nadus7WVo84UEymJCpztpNCnF2l7h8Iov7D+db+4uhDMKDoFF+4rsd7AD9O93oWi9JAgVTFh4RBX
jgRV2/sN1nGH8E2Ul5Egt5CxSiPtKgGpI9NjQbizW8UMGn3QDRe49FEXj1J4aGJbRUd/PPuVGR34
Gy5rYQotykdk9xeHVLVJE1/IbamFCSFv4nbeq0sFttktN66IjSTFgb0ADojxEDGr36Uyk5+qhvB/
8IWSjQfrLPZgmnBdm4tU0ZBQXoUY9uAgyd+307suKmbQumheXEYOCFMmxonBzspNLZc0i9837RhX
tfbp68FuOWFwhTNnseM8tZp/EHboe3wvnw2UqQ/Z+Oqv/K74saxd/gJFo+VWMnkfgIQBDxJbkaEk
6VQf+uP4N6D81px2M3PkQG+vKXEgHNO2M4WxIt0CkvbZhjASnEpLHrXzY+DuxWbOGQjHSuh7htaC
CCe4fbclsBX3YanEM4U3A0S8naDhJ+fh/g9/e79olloLQYApqtYrqOaX6zqDEHRcty6/WrHpUXk0
B4MSojysqf+wu9qnXuGajaGyGC5FufNlk6TuJF+lLCaUbG4IO3bUn5osxx8Tb+R3tQw1lYTv7oXf
Fy79+5QMDjL5HHtVrgP2g1Po8IY45d4z8UYzW++5QVIj8SwzadbjutNVGbdhTFk9Hw0o5DTOdhxM
c/nuLLgep04vDclo4Rgz/aR66atvoWvEyr4vNgOay06EU5UfxcPPmD1rI0/v3uNv/LszflshXD+A
X+WogAIyCXWr1B7bDFEwDAyWfCECMYfKUviTuGJjXQx6VE94p8G8w0glvJPl8jcAC1/rva0rsaKf
yYpB0lqq7PyR4sbPwfkOHwuDJWyNmjak7dC2Dsr2Zv3CID2M0jbBSPS3VgwTgLn0ea/YIB4Se1ns
Ccqq6eVNSvmCBab1VW0yMK+rtZ1G0ueoPRoKtl3CyivkodBiyPoXzRUb+iFC55VDH4QWE2hJKBpb
ypfCUuPLTn5ANqEvL5alDr+2NdZMf/oDhJxTgKWGBE2GFHIb2Lt1bAPKWGbiPJ4+YRB3Newh3LNY
mBHJhxcL5cRGzpbIX+0Nr3AEEZ/S/ac7DI5HZKWQjaDBtEMTxkkbtVJA0JKtzaRv8dr1pinTVuxb
KRCcKqX6qhlxL0g85EMACAV7aRhbL0HfJJ+nswNN3puYYbREihu8WcP2A3w7BsA8VpRk7RNAlEZX
P1ZPuVzYsujyKjt5dkFEP4XoqTwu1Ui3yyQJdMIrGJI0TXUnC01QnuB53mJXjWzdIEloW9POURP/
590wCCevbDTmg4wSEV3kB+t33jsw+M6NWgODepw2YyZqgCd4BjYQ8U8Lffc6acB0gZvK60rHeNf+
SkIlCJRlQStIdh2wo4+77t+Lc9zHz5m7T2YBUCMZq3W4qrQFkEc7H3JyUUXoFSoEqOsEW9LuASI/
Np5uWhcL9dl+Q8D5A0tCcVCPkmlrnMZ/L/amBBm3BvuSZvvI/af6mATemrE4uZGSSuC7tdAwL1/B
KYxxvuhXGdB83Pi9pY6wMeF6JyQFdUPKkW27WIn2U5UvCuIBRZQn2fit1s2AEbT/KkEraMuWivXw
t1sI69m5aJkorbqV9Xmxlxh7Qltkc3BX4a31ymkDNwYG93kGvlKqupBLpDt0L7YpXLpWhH1gQcCq
YruUzdkwe3PQOhrcd7E+DjMRBhhIwjA+DlufZa/NBiaFbDQMtMPorkn0ivxnwCKeY1VuJpm2Nd8C
7fEoCsbdzRIsCLMwA4gpMuSad88AWtaLqiGDK41tFRUWofdDnN8gwZhveb6Q3gOe/vqp54K3vStE
jCEwpZwZeYxE9soUzQrx/6j5CvwUI1TodMit0WVn+R8ODdKsu6EHOIYOP7YG5vJGv/utZ6AOBDJU
uwKLQaB74gtCB2q1BMyryaLjH36QLdB5+ribEOYX9UGCka05xWKfxvDU+q/y2bHkCd8wNFTanFI6
/9wS6vdql7YRFk/IDKIghCrF7/+m3sBGtXD05PoOF1NTt6OIkji3CguQsV0CXwZEzoxp+il7O+0W
eUh0RKRw6sF+0spvke/d5CquZmUAYJTl15BeuZG2sP0tM4Lc08sPTil6V3B6nnSLYArHF2huO+3p
BnpVYqZQBtMkQ0n1VwIl/8tEt+WT8SsGh7nAAbbqedJ/6wcTOwnQnnPuPo0EjmYtIdTTuRTq9f/i
AONuwfzbxIVOPVDEHxXVrlqxH1y+B1J9EmoArRCt9tV+tADkOzx+KIt7GBo+2Ci2utLdVPPxz7CM
uxIjWJtejd/O6dBjp3YrqdoWIl/ip4h+SrKQKdsq3s3PCVCunfIl+Jj+KCNc2qgZnRiwd6MmR1lX
vpHQyIC5Z1bM+l4QkUVrXbcAXwYRakE++3YG19yfEmO8CLWDtkvweOoo+TtmQjg8FwX846hV+Fs6
ovbxixi5OBuv9rf3bp7Ne3qR1LumadeL5pw5AtSk/k5fcIiPqPRGKdEiS22D/ordlU1XJhrnm19v
cxZx7vGiXwbtQVbD2qJ7I03NsaRyKG6Rhls56J6a4wf/mDdMcHR5ya3n3K7uJMzPEF85nAHithNq
Oo5/58Q9tsCYVa4qsLTXX/e6fuI16qXHvia3sDVw8McxX01Bw78B8YSSZaRzFUSoF4E4lMtmo6gD
oBuK6XV1XSFN0lDQBtaEkDOFfrGiXwOViJuteLre8PAmT+KMIsAx8ZiQ31KMfjjkwCxdJEDv6i4K
8DmMghBrP9dfQ7zkXyGvPGQIKgjw/XcV0VeGkrzT4FvJjkq9du53YiuoogaGs92rRQo2bojds5qx
nefSfHjw2KkYiXwdyvXhvPyGAWEYmVJLzi0qIPNUvr+BH4bg++/st5va8+n7Dja38NWuNPcOjsM+
F/xt0wMt/8obukERujbGI1jrEBhXC20Fk0qJmQCJNRT5kTJaI+pWZxoxNmILEBx+VCxZ38POdLg6
KR2H3+dpS/e6M6jSNx11/wRzifTzP2S/lGLjdM1EeEMFRXx8EyU0xok424eZu2Y9lx2HPyOlwXX5
NZbC972GLeN89rO7hONGvpK56MYisMeGonEBeE5v13IlZ9F5FGYEBjZVIAGcYML5xpAam8kWLTtm
Bxl9+sTA8byRw1s4BNoinVVcE6446r1HJ+lxX26o/zJGh2p6vXROeJM3Kh8fGIud8/DCvlu4Ek4P
qr8YdKslJbGt14TNAbNLpCVeuLHz60GukVQzZZnFP8IsOr+B5wHEfM2xuEmU6mbEKyfsmX2ZC8X9
vLPsFbtcperqG4K8P4aeJ0r/Y/Et2iLtl9nkHSs2cdBHVaenNaIlP+tGHztfc+qQq8SZR8FKyS/N
0MKnd5g5/klefcmS3GveE9a9hiv57ojwaczGONUGdSPqI6rgTCjJO1hkdnwVWcNeDGMdXTQ9BuPf
Hcd2+zJG9pEEqYnzUzAlBUCF0eqgIOzzQpYhWQ8rk/ziG6/pXOEtxbxXrCQkc9p3etUbyyowri6a
UTDqmIAqQh2f1KSsgUBR9tB0yCQoPLTns4/UZoOpi37VjX4apeXURI2u9G+EInpQscpVj6lm4Lh/
xDHjIsOuUDYsLtcuUa6vH+tzDq6C4yme218yYr4SyyKry39Qr8GLgWsFV2nkKnMqK8SHJ8/2+xMJ
otLpRcQuPwPMxj2Qo3cLwvcAiZfkGpYgUUh5t+6w0bF9fTYX/MLuaAk3kYRH2FvLnG29mCRd3dGP
sn5ytcoia8a2nAIO9SpcTLqcLmhvD00zk0qLCIKJt1a81H7QfwxJtfmv82B9XVPAZQIg9CaTt/+0
AjLED18mKDDp1RwfhdnZ5uNSKw13PWlOE1VVrWuwR7qHrWr5CAKwlncGu/IjqWb1I055Vk6R2rDf
iuyh92lAMBC/0+8rslNU2LjrhaxKbq6paOHyCBQ6Ji2vuSQsJ1GTSiyaQdZGTu5f/hzcyMqomB3d
bYTZr8o+rl1qXB0Jb9pDM1lrkWnS/8jTSEN2UXC4gASOe/XPc2ilZf7sBUg3d+sIRT/3i3gwrE0B
J/hAu8vXnLyWfq54nJ3sX9JJFlswLOuzuyU2YCqYbPrpzjRi3XQ/HD5/FtPgbu5sSZqhymMmkK4q
XRmI+DIMV7jlr0ZRLkhuOgrHjCc7BiImcIAJvgFbCvNYGR4Jw/OwFpNfh0upilcrXF+wu1CAXtAs
PLmtgn/g/id9AV6UStAdiWNQQ4XQOXONxo4N6rKM/0OrNUFac6NICOlchyjGX6qJ6uIVh8kXTbOX
hUZ0JFeiMGtJI5pI1uhDqlR144b978pe3zIzjRvPEa8qOq0n0xLwCDiFUZeTl54MOIFHL8T9q+Zc
dcXS0VaDz4HbRZhumA3cC4EQXbdTwsXwQD+kVuTYBz9eeIoCzDa4DvkM1TA1IBflNMpRpnP+8WaK
4jGM5fDKjvWHJRce5lmVjtFiYskEDCJQ5hnmgBGIbMoMs5JhgikqaHqhvF+zWEs+/vnilXydZ/BW
+22/aVXAzYRpcFkLI29wtvT5RRPIVSfUwDAdbHex/y8BevvEe4W+cfmDaLRTrfP+i4Ye7yjJFD24
xsWdViycvcCC830Ov4/Ge+8tBrlxlevCNTtD0ATTHO7266pRIU2ogzWbaIOTtzfwZUBVTF/XAVA+
kHJPkgkKRCcgc+o7mSFbEvaj8bsQ9mRO4F/D4h6uIQuhdkLlLh4YKKBDOVsIR/Q8wR3012IOiRi0
SKpvLm6JN96XP9Z5jlFs8rAdx4AOlG46wmu6pEI0UwatAVX1WLgdcqPZLzo/v6nmm4nkqqQ8bCKN
pnmdV7tUm1mPFuOXdLsBmApM3CdJyQ7VHWsIExatTWfeneqXMMOZfaV+peuA6lhSkz6HtYz4JpHE
aQd/DTM/D4LbHYkHxlcF/t0Z4bTsal0GhbyrEd/tjIgFv9bYR+1cDalAt07DHFy8DF3tC2NSB8c1
pqP0ry1LJdffK152ff1kZb9+2YuXy9bqgA0KhLMEJHo360ez+TFz4DkHVeCozvTQB+UozIrjPgH3
XVPxbUX6+VWD/3VJWJGgtc7o1nPxPzWicAbGIxi9FJqIzTlT5WlyaukcuejbIraKH23h+7OE9gfh
aU4h5xAnJNp9oR1/hDxbj3p0qQ96eDRA3LvaggFfNj6Q3Y8ZqAwWXBlt2vFQezSFidI9AShIoPOs
cDsA/SnPRYDVkSPhDxfCy/gprSvT1Ha4DgXR1NFLv9VCsKw/URBaSlD+ADanHwVAqtbFvWLajhtn
tIX7eOMfclWtbFfkRXYWpiWqyNkpIxnsBeY3kRzeoo/Y5HI9rVpp9FmoSse8A8CXsGirkSZP3YwI
OmdR7SNF2T4fNVGlUwp9rGHlj3Ld1Nxbl+IjuzKCpi1NT2Q2inrW/7sEZIfZZdbvZJs6UM7BrX+d
+i53Ocx62EMdDKsLbsz0Sy6zZS6SRAWIMYs5LPvybMRE3zjKqgJah79Afqyu5aRLvQ6CRg5DMu5X
Wtzx/7XD5TR1fRknaRVaq43LG8bigj2HwEBuK4JcMmA8E+tInDj9zhvVgAQ+/lOwRqKxt7eGgBP2
DuxprnFHIGQAWP4A+0PHROXOoQGK2uvm3mHukmq00tdJswcCl+ZqpGrLaXe9aA3j11UfmshLXUA6
dnqEigzyTCtybLKT+gLWFCziNBpfmUoW3tnCeZoj3o8QUbzTfEVFaQ0fjrfld+oTm5m3u8K5lKYL
PqM1K1vepMKVdWoYGJCV3Z8d4itYc7iBpBR3H7fuBTukwM4ck0c34JX0WZqcgxmDGKD78PNyK9i7
0bav671mwQpbWF8BYcWWXXQRboODC69Oa2DGImMFKj6tl2gA/OSqBWKGtlTtEsaY3SksOepQYMC7
WgepLCYgpjxnW6lFaG5UNsUW7ezopq2fL3S+Zyco6HqRMK5SmuJAKiF9F8/U032qNs7yG9XHKv3R
luQPVkfjL6NkADCLk5GPWUKT/agDXVNKDcCa7lC/RDqa9aXQskjr/tWZP3+2UCLW5XyLCFneR2JQ
Ymny5REHgIobgA6KFegDm8llrSx2pMxJCFb8u9rgsJDz8TDFnOxddDcztD5y/1diYKg7MIgqU94H
tyHkqSw0ap9AWhO7ybfQgeyLM+3UVtA3HJXapWJkgsWAwaoHDbALrjkPDnHPqkb9Z+8xzNzrj1TH
Ff3sEH2ZkpAachWX+ZuEJkToZY6i7gy+wtQlj3F2SdM5wFRmMcvWnhNVMQ/s388hi1ZXljmmMDnq
he/dFewMDxJAJbl1F2jWSqwBGSnodUCFiOGNannqe85ufqVsHlWSzdbMqJFulOFg/3kMAKdPXI9+
xOsSEG/BNz1LmgbuqA3jLWJyQ5M5FYEX1SPeBTEywxS3C9No1Xjy0211A0KUsPVrPmqlb619QFJj
7L2zdoZSFFjHZmIsLqiZo4C8aRlQnnSDhIOr+EeFut9BaZm/Z1AfZJsA/RRhLQlxTbHr3Iue8OBh
SDceZZ6MiQ/a1iIqy4nI2cizq5AqV2dlrDjccovyUwTc3d2M1AER+AOvE8MivByMiKasmz2vQZlV
Q4R0HMgEYl9Xi0y+rlgO8gSld68LMHrQU16BkJg1zI7y9iqqW8WX6nKtyPIGDUnpJzK0a/oyLrb+
cy0azyZDxtuwGyBYeTo0abcwDjX9uBaWeT4xPF/QdHKyrv1Hnr0NKRBIiMmufpPJSPOD7kimrLkl
lHahhWF+yIItZGbGXS+OWFGlOIgfhAWn4/BMxXHbh7w0VYqEh9np/OyNHZz65TUzDupBn/kiG5zK
CgTGe6vJjBrny78pxmjk8t4i1wOmKrbejObytb+sMyKAzDDwnrNYspGXRucB4h6X9l0jxJjxhTvC
7B6s1pZ9VbqUIen0sWDjJL0FyMb8wzIqJiRi6Qz2qqGl8fL9WB8+F4P1hILqaQfGmp8+6gVGmqe5
XmzjlNWMm4htx8MQR+6+bYcAxmCMM10dNn8qwKASXb8BrQuWnVZTve50YvR/gxLMVMIa9HP1WJIi
Q67uxqy41LVYUzgUkIuKx8m0SFoBfwoqNJUqE4TH/OVPy0IATIhFInW6ZizjcBiMAi7w76py6Y0z
VshBBFlZDPL5szpMcjPbTOyqE1Oo7B7Ym4EvzNKIYi41UNwxre7TuDkvYCiUNDlXSDbZk66QgSRK
MsxKscvZ0v00V05Mrb1M8bKBCE7LDU6MVjfqBnCThGQlI4RR+q/9xkYTtJgXbFZcepP+BzVZ9qVC
899yjLVOP0euYyBfXzaJlUi3jCYu69ovckAynrC4wFxwh71jKxpeh46cN8S40/TKc/DmHr41bJfW
jqY+Pd39lLVF+YMEHmDMy9mFZfg64as8/CGMLiNSboQPCW/L8QJxnqC0oZri8x8lHLOS76gTzDvE
i/34seaHVBjGq+geGd7K86gbO45S0DjPzDtknGpFNe4rTHw4Oi5ZOu0bO/TSazKze4+WTMUIaOTn
jByv7s7xgCGGSukth6N8xNZiD/sUcveWB9zKi33mc+3Y6rk/ykkvEYCK/ACmFtG0orO26+9CrO58
qp2tf8xLCCWurz66MeXZPjxFNrLQWFmAYDPMVoXAPzRQjCnCZKOcD6UCnKUljiVcxgxXCwInrPyR
V9A3TQPPYBX/J1GkMHKycKllzDHOmJbZpGxXIS9To3KdWe6lsDABPXqwx40G7SG4DKdgkPNOvDnu
tCwmBII0EGp+40re19p45A1uJFK+363FDUjz/Hhw+dQYcdc6x3iXew7aKOX3J/W5Lu1wIThP09jW
SJES0tVyf0h5C/UJ0oBWFD3zu/ohOLpB9CKLqbFWcTm9F0h4spXSKqty4g8Hdmyd0nS2t9mhrQZz
bltm2CX82lan9O9ujQhawHld1eS5wb57EV+og0Czu+hw4vz9YaELVWn/rXAGahwbUeJVM1tK/M3g
roNLg/YAzwGhbNsvbCukV9+xChUVTfxkRtkpX6RFFfODV6fnA1zeM4S15KGKTCGVneX4J3EOnw/r
68G3c5TXThsYW0U4jnTmCyX/b/bMK8qmEcjpOjVJHz3Y0WMe4LOT3VTDNfgs1ruYBod0Ec4nYo0d
gaoMJvaWiYj9oIAe3l0nApPQin7hiwbY92YORabOjOSdTHUxzQvLKQ0Xr3JTWY/AYZJGNk/raqgB
TNM23WfHNnmrxZ8M1QUHamMZlenIyrY+O9X9BcrLLyNVLre/ieiZDiBZiteVguu28nGzZVtPtwbB
457OK5k88lE735KIFBeMDTPiX59MCuDuHDgNSYJiKXjjPWLgbubNGfgKf8gqoM/fdlkLWohaWjZV
aZQUiQ2fk6o5O+wF1vNIjTxKosWtNpHsRnCYk2GywcIYjqww4CxzV3bpCoJaphk6LDs/X9Mh7Y+G
81PFZ59wcHj/lK5wzrSexAJG9F2o963n2gPat6AlaftKnm8YoGStA32BQjeXD+Wl7QbFIgzMcXoL
EXbnOVbJEMcPE19TXNUUmW2ZCGFLLMaBP25mHEMXFtigOO/FEF0FzNRbdIPo5H81kgMXv2lobNHr
vKaxSVZvMEH0eaMk4L078/ndlwbuFuwBVCDkU+7NbD0F61D8JhD87pLjJJpelOJVQVPPoLr4tkeR
KsPnQu1rxKboT47QdOVnnMvP+uKB1xKGGmOdTHkHLllC7Z4Vf2qLngiqxsWmdsQ/L+8RFsW3GGdH
npdNDk/HuujVQc2jNbQ/ckXU5wKH28oarD52Te0xmZaITvF3vWXC6nblOCODUQBQMGaoqxEcqXUQ
B03y4TFuwdOPnj4XbXppAcYYxydty7G9pgGA9qw0/WdAKfcRb2VeB7SrlzSV6xCxQ9ztsR6bxouM
YmUtEBr+mvk8G/pQYB5hmdGImd/CFTArmJLKkTu5HpET3YY1dOM+68hXI5KfRNy/al+jqW9v5nI/
K5EIxgx369PI/+Dk+5haVvZBGm1cMLjawdx3i9rOeW9vOE637Y/qGSeqnWOwkxr6H4NqBTQVWdez
eAd3ekRhC+1UE93tLCkhFueYJEq15wtac4du6YMw24j0ZPyz2iCcsqfV1vku181aj5IhHRci25QJ
VB1bv+mn+xNSGHtHjTtvJb6Se3BCGKTig8GoA0x5d5fNxKNVSIQ1ExWx9kUXlhBLuewviv7MRVnK
+E4LMf5UFJmh4z2Ejzna6b9W9KnZN1QC4qIMMe8wfu0kGjrALyb+IxPeq+mAW/HA0DyHLqv2J/vq
UAV+xkZHa40CyeQMexABVXGSCwJD+f0bO8RX3UYA52SNwVql0waP3O9jovHzzAwTFl2soacOdXJf
Lu6KN9NgUNEcQl6LenyaoTwBHtWRvK4I3zh4zv7LYQFlfo02e82fwHHiXrxjvUwyQ90ZNa2xY2nz
h63gpY3S+AudqZSeYN8fVjG4j+TorgFoTXcaEJnB1HZo7EbBqPYxlU3P0JKkuyzg1nWvQ1RhKzOO
x6JPITuB8otuWt//e5Bne7i7cujFzZ8+0g0ZC1m0LJKlZmyN7wxUalzd4qIpOTpxsaTAifKM4sOa
LVYvNpdmG5pjheXh11TsavATsO9DaZhDJX9wd9pRicXuxS+gW25l/8+ccbmBVBqClMFrUw5dYOAg
rLOStnAwX5it8ZuA13YP4grRirfYFe4W533DgQHwx0NHIglZWhHrJD3H5tWo35qyCyl5pKXslVnb
rxJu3jaDUa2qMjBQ1EWU1A7rpxQM/JKWCdrk5VJrjxU+DrDpUzkk18xTrY7zSyuuaIU/fyZXbphZ
ikRZpYM/ZSk2lPitLrEelqLyQR8yFbs/rjmQM2u8Ns+TI2YZ5PS5yG9+4KX2eVtsUD82diHDMGrG
bnJaNw++YGDWmsEXKSWdCdE3utbHtJeR3qv35BR2cQI628FPuOzFei2j8yMEOA+ZxPuUIDyFxd1N
7jQgRYu6ZMeA0Lb3DLd2E/GXH5/OZGTGjstXfuUtfozWM+onEsE0+e2P0Qru8oHcVJNlRzk9MNyx
/2uRuPsVgfQ8gl+Ra1H/b2egTC6FtlGfWlitBI8S1QLLDsysl3nd+Rauvb+KmaeggdzFF5OVigJ8
g99PPlolK+XUgYueiymRCMiuSNx1pp4JLH7U5LetWehzMrifSSM82gSHxJTiWThGGmEZsm6GyWta
XgsSkKE7p9j04HOi+aD29bk+EFhUifK7JGO2cmUXXfJiT2+7+Xi8RdrgS4Wcqx7MMrkF65NDHK+M
yK2DW4coftL9hzUHdzNFog0CH9YE2yFCm47fwM7xx414nC9wFnO9a3Zj72D7arHOKbtOmqqf5oML
9ECZjP5a5QQPGOJOd5KeJPkzGz/QibcXFgt5FR2GdrXaymYQbyhNKDQyLNxYIqcuLyfLD3/CL95t
Cl6S7WuZtSSIjI2lGbLAnMojBV5Tyuup5LgNjrNG08sPp13PXcj15ojC7V5Pju17W/BJDbBHsuuG
w3oteQBdxOq+7af7v1ZDDnVHCG6n7w0yWyocqWV5vAfBPy1aFjgzdqD0k6ixH6dKFe1Y64vkrwW3
Nq2N9hG10Osp5zAnITxjm9K7bm5p/0iq/f/CexIpjf1lAazxy/I6KjXKMoBG4p2UnhynT+z1VQI6
DXD2TGmtwCfCrjJwkCepUSDQq2g/Smus96X0wCAxwc7uXahnz7vtEt6hQ9AwY6+3q9XCQyKAJwtQ
GIww7U5Wy+saPJUMWpt2mNhiZWOO6GkKg9QWR4+0jYFT6jKlUogTuZYGF6S/TIgqBMv7llLMaKty
0/ElrHfE/fIw3nWPTftiL285pgTsRCxsTTPv6OpXVFkFMbxfHtCUMOzYrPfNSN+qgLYecqwsuFws
SvPGwfxs+v9jnbnk1CDR/YPTRd1WfXZOeiq400iPudU6gNHx+lfyFz0pOKtcRjVoOgt97SnR8EFh
cFgBVgikXVMXXfX1svl7O44cf5OV3ThpTlmvpksHZRNfdBVQo7Z5jF30SRJX7ttqow9FHE+azp2O
KInvuCQ6elogHooh6ARBEnc5aQY99C09eJPUnSJIgqEvn0xsi3dqOKRx8UzV1UC0wL2jxgLjeLMe
IsZp32XYr+dzEFSs0ABpt/uXSeMwJkjzjAOY5Wme03wgSsWgg5dGLV1Wimj0IDm/87FaJkJU+I8t
nDyGrBef5KQm5JLoTFz4XOyxxIuL7s4NEk71T8DhD+THHuXjrWv3rirvERT+nA/Pricdi4lrIBmK
xwM7JpAeoFZHtXqV8WlWaUHqgpZasU+FtuiDNpbG5qEKhHPzAQPDRWGk8ACjUEUpxbFlCY67r0aA
svo0NUOJFOpdNIZv1huM21+kicqjXNhPNCa54CcaRYiftxr9m+Y39x4B1fmzl3kddEK56WJsnPhw
ND/SGbqJrE39r71FC6XBRrZ+4Yzz1NRdvQaP3Sh9HPb9wZp9XSITKUDIuvAVLNp1AtbR7ZzhbkzQ
uJyS7bIA/AGG63MDZ+Oa2O3s/3NWlZ26fqpjFSrj6PtHV5AdHsal+mP1LJghq0h2qUE8xDRYARmn
9ero4NtD4gLiX/J9TQ5MP1I1S9XHv42oSz3/bissB9Cm0ALxDHhEwJzNhC/nacfy/OCJLxeJqGjN
/+QR+J6XwxQEvMvWXkRh3M5cJB2VGL9WI9THv+JIFUJFcJmHwi5LNjhovb3oroDBR818sA/keWtz
nHCor/ZAAJnmS1wVYpU74+orb54J8TJSu6mP7/6ZP7gSOtPxowXDojbVZgcRHts3I4dcubUKDdEe
y3L8hTJMLbPMBkB+rIQwDzSaQ7zSDri3kJMcyeLzIcfyfFXU58kkt/qCsDn80qJHKJ15E1v2a/+W
gKYVr+ooCV2w1yof/3JXlDR8DrZvrlwkVmIaaJoKKr9zGxT5jGaerioWIPB7lcJP3PAKFIPaq9AM
VIcdnMzPqPTmfF6hwc3GjD1by9wCCTPnTBm31rmnK3F6o78qeNCeZh+dQ+b8MBXX+MTrJQLDPIrA
ZQzS2bKYvjXPPrQpDD0gW1IQylMMfg2kJwPgn+gYDxXNmpF+oLjQZm6n1K4XMiU+n3vXU/DH3sGr
u0AJ4E5xY0A1VY6kdTpBO05copPG7kwuvm9cIxC3d14HEo+QJdMii6behxkvDhJUhqBlxA/P5H8q
zlvmEVDBx5ZOspTSTFHtI7Ks4JGHWl1QsDO6aQa3HgPPgWwMXR8hoR7NwZ37k47n+CRk0ovfKOzd
nx3qJiSjXkZg4AC1pp7lPQgkVbPBG+8Az2K4qQ5S0B/pi/CPpLZQCAE7Eh2OEtHeyXNS9XMcisE3
XFiSeThn2PrZeSXC9LEAfj6XXpEZJFRR36KvXDOL6ygMSGG8myAXXuK4zkLDsgVsS2l7E393YUzP
yZe4lgWgkQpsqyNBZmIex6DsSpf6Lam1ZXKqiP7xejca+neW+bWwMSW7sAjQJmEVENrjQQNO6pwN
nlIqpdWMsAtMcLScwzD+bSUEENSGUSEAGLjy4uKCWoTWcLgQxzAdlr7FcI8RY8MQ2Zdx3dMuSS87
0ggnbkFM3nDqGEuqWPkN3lkc/cO744MHSoubgW4/8umYZrsJaJ+cv63FyqER1dHKVcfIWGShyFBa
0mgUXT95hQ1lcHks8U28CTrDiXdRPTA0wNDgD0rNCZtWdnlVB1yIV1OLlVYUVbYrUCQWyadiDZtd
tHtis/4Pov8NJf9qJ187lB6fp4mz8Gydqrn7YzB9m18Crc4EK2l9C4JO0v/84bqjX0FubTyM/S+k
T8GKJxk8Rk0qkFYQZ8p/TyeMZ85SzQRNfvfQ/wpaQON37gY4HQX4cY5Lm05wk+aZYvhsG4yI7Yuj
C6XJeaE3GOj6n/lrmC/mxxEzF2lBpm0hB5JeJxhvz3XHg3WMcQVe02NpNJU8ldOyokAcMi3zEnaE
es/6Ped+jUl/SMp8776h9UEigS7P4EQg80TBtVNUgUuQXVTCQCk63ATeu1lN6hAnygWrLkjEC1jC
oP+Qsxxs+0iGASukwll7XBMgo4uNYPtiY8zdy4JnrcMBF/alBvMLW6Sa4ZQzSoQZwDlLvZEEuHsF
q4nD5VqA4Qha1kYy+KE5T0VbMkJJ5wVRmRkIWOlPndbPleVSxNx4+/NDtJG1j21y7/vcU+q8+JCn
ngkYHEDCo+ZlqvlY7R3h4S4MeaJvx7gbRFSLWhnateafBOBPzVn57LiJWr/jSI0Xa8/4VjUCDZ94
yPJpbtFz0tncCxYwchF1yUEgCCxZlWyhg5tNbTm4RG2DwhkNQmC3wakGy4a7eRd0hXiOkXkXTKyJ
Pzrl9mdoW2QaR6+tbOxovIDGqkcIy9/gg0DpGEGKRvIvRGoig3eoPc1rHTrAzGLYb8YZOha6Ta8R
KWqR2wuFly/kHUlIZve8/2qoyp2w8lldQbpFR5LwWkjaJ/QsGTYbW4KmEZx5Umm79WD7m/NECppi
nd/mAS+e5buw1SvYX1X5GCsaPdl+gI8iU1MJNzB9oVnEDbddvAU3N8wuO57tgyGuCDE9vwhNz1uM
dKk5sqheTrSqX4WwXWaJOmITR5VrnKDmUt/Ez6+EQDbDIX17ms7L3GjfD9sv5/r6OC/CPmLgLg9F
XGasnMl0ye7I4EHr1Ug6mneoU6MdGnZi9S5GuYnd41VntnQL1r12kCI5dVbSuxe11DbcgeBwFu33
Jup0SwSQoWUwfh8IBQkOUNK3TecXr1ARd2a9cB6MHDwabzb2onOvSk7htG3+qhkkE1i6zK85nnmB
+kjqgjQNsl/9HceLWz858bSTWnScNqu5hM9PV6wBdJWwGlOWFaXeDD2NGSADzM3rpGhctnhCKVOe
rHakX9/nmaxOmPUC04QrE8LQaCwPRciqLauqfF4LgHFoxCF06OUYvyDsxUbkTu6Jq3Ren1vAORfI
Sn2tiSPDIffeJ6hNBuKf6VVvw6UGiXTT++GQ9Xcz5omoHnCJknd3ccENuKWWkg8YujMq2jcfSsR8
EwhlVnP1rOnAV7aViBFvH0aqPTLRFkel1qBgSyz2ZwkINlSU5lLlEJmF1ehCzdx3q8TPY1MldZeg
Qrn4KHEXxB+CfonV3/+bmXjTblwCg1ewn7gUQ54L3HTX2srQuaU8yOds1n4wg2ROZCmxo7V3JRYE
e8Yx39NhbLXmXL7tofA+eMdaXRhldIWleyXm3eqENl2VpoZyhd79ZQ9UPaV8nQ+EMhjAPLB0cevr
8bezJmBIV7rkejWFJyzNsiktrnmncsVxIKmuCkhBXUwmqolBxbU+4tOrdfPV5s7pPpAPKb4EH7Ks
+L40EJUQK8GuS9eTkVeIoX8XIrh/E84IPJiFfi60u2V5E7CdiEK8s/neGl5iI6dQ/ZHyBcL2Xksg
9yVLnVLxYqEbLTHIvPjl91YcBwAwPOHbdilNyTzcjkYwiwMVJx2Ns2AB9TKwv35Zlc9E22P5H0tk
MJZuUs1hbuJ/ICBwFngMHWtao9yp/uiUmzJvRiXMcST4AW17iQwmWrlU6Mm+IY6+J9/gdhml2qrS
nb52fISxY+BQRtiKkItspYtFfeGp9FmFXD23Uu6ggsHhyxmY9KC5P7mFi/9O4wiaGRGwc1c3MtOB
ID2MsYUT6rVhTNGVHBX27b1eix9zx5GGhfM5n/k4f+8JZR52D3WFs6PYzdqpx9xyPkMuXk/83CCE
ira6+kzPc+EKIddLd5vX/ygXECzbJRhZXMDYKYiPHDKC7KRR2s4DIHwjwLzaNodM9mEH6iRVjgSC
MbgiJyTNNQ1jv6JEu4FjFZjb0wYcIBf/vDgAT9i/aPW4Kj8z4MTrN+fLL8PzLNdvrmW+RPZGSYF7
W5+IAXoJDEMf2j4tawwljWK9Bvdf+9zPcM8W4deD5R4ewjHxxOO4vKiP8dMENsVHTgmG01rVZg/x
2OccilvKVuQvLhnWiOZuWCBSYEiYTxI5HOU8UJ0qwfgMX5vx8Hfzz6LH9QK7zDzSFcCO4hRHFHcP
t9oaznYJiuXYYgNqkdM+0c9z7cf94rVvEdlEAJPifLk9QwLbZD/JasysvcOibJiqytjZBqiTqRkO
2/bTHM5VZ/wGQpZpWpUa+mGYxYx43or9nrcdrGooTOi7fgOUdViLHIouq1lebCewsSPftEGcxbzd
njhNLlw5ufrgNiEEqz4EdDq/LieMwUe8csAol67QPFfLdvyy68TjP2/qWkfeoYXrK8YbltVtG5tM
YwnNhbUcis3IxDTvBzf2tfN/JXzryer8bhw8w6UpOEUaFTv7cQjwIpp01qiNfxuLhP72TPCjXbbR
nK7Qx7x8FYbR+LYrbPXu/pu+1oEYqNN2surFVOtnTWpbPDo6Oa4x8WUv/D3P8ZQgnS+nYQ0GKm4A
MQNbG1Ph1r2VXFCZ6yHK7hcWW1v27VFZ7m6FQm9EckM1KToXpq8YeZF7UzHc4wVTOCph2X/TKPg5
hgUVruhRHoA+uBdaweWsazRz5m38usv/9yN51p8o4DJauZUeBtDlFxiZuGV8M46bhFzw82XimSWA
JcQU01jVDHa9Nssu/wDmEykjeHh0W5d91sH+HcJUlS5QZODQPC1LyV0v6SolqDM/6mvqi7A6EHyN
Q4+qvQY/OAdhEe585Cn04wqWlBtYwhWBvGyrEnPMtwQ+K65tRQ6Yij/rs1gKZCtA2RQlon7Z6jSe
0PmOs2D/KN5plv9IC6rn8QY7puHMqlNot9e2XxRGHtX0bLBavSNvz3G3Lg83ATSWEd4lZRFsEU8U
vkYuWKMLQyGF+xHHgYQgkDI1KyNu+iyVBqNVLJxZuw9c2/2y2e3mo8oppi9yZd6WVat3utFsj8Jk
EM1UMSS5y/5mT9zhruUHZRhcL+4O0I4j2cN50ZPSUqaaUraKvWTVTdqcNX0BCSTmf9p7RYXPgmSO
Mr7M5JVsxZroxEmNb6vySH2fMesBzTaXhMtWUNnNMOQH6rDXXZSYvrZY7PKjqj0NBWXdYf3hxeuK
B8xCCPuk5GBDbtsBG6y7jhBX1QXjphEnCHQCkCJ0aE0t5mdE2AXr+Ud7gDhGhMTQPOoF4a4W8Idr
8lV5tYUInnpaqI6ElUukne8I15om/kFSEUuhE5F8tucyMpgmQTk19JYjK8lln3h9nF5e0Ex9X9Rv
YcrMCodQHML2uXM0gScc+ZFmNsNgJVEEiJ/XR71Id8I5Q1Z10RVSrx0+IE9PWDDzAfuzT8mOcunl
uy4eU16oqkpEZ+GIMN0QGfVF/jP/X6srzQepNPJH/O9raYVEaLKdy5y75FZ9Glo5S0GFZbkR4egh
Od8umvx+zhb0Z0V8Ze17s4vwvOjtkJLTVI8CUIhWfoPszXbzoBkwuwecXmgTi323VKHD7Y/p0dxa
w8ASWGSUFzbofcFaXE3mhl+MAlLumT8SUaxWmQRVZoh0irESpSgEfcaXUe9qC4SiDLMd4a1Q9P4A
YsZTkNjwLHG18RLHAVGCN+Wuo4OlXbTesv/A9KRkdqFe/2M5KJbV1khaeNP9CW7EniV3q6j2km0v
c5ulZm+BDQGccORYq589bdv7s6PWd50xbhNbcuNWK5wLELmSDGnBfC87eloqcMFVOTm5SV6lf8Cm
zaat1UfAtOJkzEGoWBK8a+P8tbhnxD1vur0/sJ0zUU/Yr1ZQrxrMqbruCm9h+iszjV+PmyE0Z67s
j+IaPu6xM6QB8dT0XBS97TqVCYJc0OKhUVm/pE7VtLlBs6q4Y2+q1uts/TkBWsxB+9N85bsaA0KN
Dm57xJ+pOZ64FKA8NpgForiULRNNP5dOa/YwryHaHNrmicpzvEjMfUwaRoCNYdLa/d5iyXywtzUk
ffYUiC9M2smrmhlPQPml+CARWD6xY08FBV+uPydaCeGkUZVWdfmMeBjnWPfD6PY5aP2bCYB2m7wR
3zSK/Y/BXJIg0Xizk2O8Om86N73uBHFO/QC+4okFcp4dWuyJLcGt9Zg+crAccp0esfUXWLVZTX9L
LuVPpJ3s9MLE6Hfr3uik+LHAsRvDCxc031UPQw6nzGNz3RppE35CwB/JA9toQnt6ySR/BP/sgmYs
Tj4zLrPTF+L9qwrClX+Cwiju53tR485YzXNW0WqK4puTqUqvwbjd56z6k3UyBM9GogRFY8g80Ff7
MMP4TKKQLxw3FpHKtjzB2pgAZ2WTkBygwBjkgf6lODbpWuAI4ixKXdlgeXsGJq+HYhmLqwT08V5a
1um8QdJd+2Q2rbfHy1yYeVNCp6OT71N9BH+UJ2urIMAeQ89ggdDSY442Vnp6yHgsxE4k9wBISglb
5eN5V5X2FmFCA8trfs7rRefQzZo1qo3w0qzhOM0HtsNo5bCdBzhqRQyOIMI06OjHaDv2yGk3LknW
7rYMgaK04+FHQhWh03aBsjUR7x6Jdf2kAblWTZDUiHQb7TUJBCB+rQFCAM/WYqqzRL3zoiBaj4Dj
NzJQ4un7f3hOOq045q2EBvBFLGYlHqLuGmjOzc95r6cTIUuSc0NiD4cDnOHCuUcAO/xrA2+jKbxu
GQSp7Zx+dBByjlXaetLHcJFAiYW+/a/FR6nJMBFbMhhm0KZ+8rwLZc0y/W1AUWTsVFiQ6+zEheKu
6eHRs3VP/N6oNIJrrPzWN6CBPBelyJofnCSodP0G/43plUSMNASDxesOQCzBX3a8X0pZ2aCFe/cI
9SJFF7kSu1jRglnuQJnRdt9d4O4XjKbMQ2XguprCcKUfNVNGbgwr0enEryoWcT6RIHBKircQjqnT
hDR1OogihQ2aiXj77RBbDJa2l+WUTxQjQR3P966NvCSW96swv20MK5GhU/+TRgsFtsyRvejGTTbj
jB0L3BsfL/Usstd9N9jZnXwzGyNJbZrdttGH7t+p+vJElLio3pgt05zzM9FfF5PBqN9wTNXivQGb
HZckvK0yZlWtQnJJuT7ccrkIvwjpTS4agznLb2kbmZFCnqw6qRriQ5vYBQEMOlHzYHAwppc/bt+r
8CH9aTxssK6IbZyAXIUo9+0HPdcKz8rpwLrXEgM6+DPU2JZaBUbsiaRMGvr0NQdkqXoLTzTbAkJw
3wqSTFhja40YvgJTKctpEdMvkgRGc1bzr4QFXyeg8iGAIGR77COa1rSfx8FEMLEtg1lwF57eHa1S
gqkGW2bm6tscf1o+rOlPZGoV5Jl4d3TJbKc3A3zyOAzgoGeuGCzDPC4LncKEjroe38ElX4zjZdS1
7cACuznAli1FLY7JX0nAiavvgU8IfVSeN2h5kFBT29TFvGdMDyPN9lQDFeIssoH5aAHnFCnKGbcU
EW6b/iJ5PXrHmrJFCk7lwMEzV6ZP/sbGnYeTmvo8/fT+O9tjCPUgDKXwf2/hwNPHjWOZp6YyQoXR
LNGD+tJ1zV069dGthDAebhn20ERFaw6Vs8fDtJDb0n7Y6g/nZxp9Q/Yf9Jji6prUHxwBQmu0LczN
jm9OZh32c8kN5QG1RJAYQgEYNocQrDadQt5LrykUgL/Uw5qgiPEs9dOT8iDsA8eBBXThfUAyPElJ
fmklJlJBt69dE+4QyHpx4Ort3XVpGHioKoOuDuHI51MkkAvr8NUv5ao4rE3BoVYQZhRBxY9jdPcZ
yU8gbQnawtpMoJVg6jyRyP47WiVjd1x1SO8nuVic+5Gosswnhivu8sVBQTJK5w5iTPgHovksi41d
9Mp/slZHjRPe2ErRk666carvo9pKAd0A9NgO94t5368QkHL0oGsTVq1gsVq+APGQc80R92mmFsfo
VklHzFIdZdPdGGI8F5Zsho5vHWoP4I41T2J1ppfMyX/0P01xm0XMZ8iCwj9/cMnFZYfxkhrvgdNM
Lhq9BJx0J47CukIAneasPgLKRLV5aKqc2h3QKw4SKDKq4niWQbkolebwIXbPTKB5FZgGzsvQ/+pp
t24ZwEXWlw4OIFtuU5ZxFpdTjUrTZYGlr0eFerLZIAQUB1yqI2VNtksvKrEud9vmxEyN1N1KQeJ2
90gxZwKmY2sDoqJVlhm/2FK9KcUOoRW1DHKgenWRV8V+uMcom9rQek1B1+7QRNG6p9Fr1CtO3W42
qN1Wtq3dxAG9KbaoXIY3mWoGbvvGHARwXmq/ybUJoNKv8bs8aACsIhGdoLQJAQnMOR9OHfUPmxsj
0sefNv8BBAMT509nAt17WbFU5XBfb0+VyR/usznx58KwVqXlv/KSpk2DJ98iwk6RUjq6KCmZnBlI
L0CP7c5OgnZKrOBCyZ36RbjcEuSWHj9grEka69LdKr+Q1h7z5T7MGfDNheLXqYYUO2Bp5BeNHSNr
KibC6fZbDRGnMtn9ttza0e2CvTgjbF1q987YE5jc2xy+DIggD7d74QPiYYRalwiMJ3brilY8eWpS
wbPOPRPNN0H8iWAIxaEXJ5mMUnaTHSfy3TmZc2hZhn/UzivCoY4I1w7/PcVuaNP3vJPAOyvg+jqA
6TGHeOlJ/9V9/ilKPUnWz5BE8O53gzS2YoxWEzg1ytOf+VsIGC/1vrFmUJgeMZqxovI/HFl6/cu6
k+5iK5s2WLB49HU06TQIildchdbNv6gOItE7+KEl0yLoqGIeZdzttah5Lu/Qf6xXyx17NYRTBpml
9V/35DSDM/SSHNdy6HvQAHuG2dTIzi1mRZuqVe+eahIO7c5r4T+8nnno3KWmVV2gbWlSKCwZ3mFH
mFYnjoD/Wg6i3DOjUZ7ge0skTAAjY08kbWW+Z8dPLXkIvzXYqR0BCkVLiGm6zxnQpPvQ5iUUSAwX
A60l8aa3q0V/wpmcFBC/HxGNpNb02iCpBJo6w395Ufo4IbV0Wgnp3i5ojzoH2wVcHL/VAj4loReu
tcCn9prwkhbFn3OuUQK7NJPwboxy9RM/ohQqGxuO2DiGlbE1OHGmEOBEeIlvxQl7+aZ4jWq3h1Gd
e+RXaoDL4PpZgpLIVJo7H37lwd0RzncElhg6tasBjHYUQYwNay+1amRcFngxzuIB1LxecGWxmVOv
H+7c7zkft+/uSmr9nXMFHMdaHdV+v2/yTKQ2VXhtKNoViMvRYqWcLInxA+2of95me70aZa9B+Z69
8S95ZzaSYeg+lNHCihum2ffyhEd9kijUFfvq5GSv5OMuxOIXEc2buxBo7833K2tlTPzJMd/B4+7m
YLuxqk63S8Z6PamfdhpDBopCUT6fVgWoSQtDhoodlBCbcXfBmQcxuRoSfeZ4ZdgGIz6kvU4gVmlN
Lg89TSa9VQLWbUPv/jgDf0u3n0Pzf9LSt2nY+6sqTEwULfrriaZuULzCkMMLtUm4kV54w6xY/9ZS
kcjQOmb2xAhoMIx12+FZLaQE7Y9x3PnoYh6ESu3UdialIS6xIJ7NGbJa4goUho04OCCyJd/wxElg
HfvYs6qFar9fRWzEYvMx/3nDufERO95qO46fHDISN/IbLhogIa07fzvrYkRrTod9OEiHTxwZNpN2
asWngJoINQPhJyJOm6m4XRQo6+koXA3KFhse6w0XfFEKZFs08oeeDfWIpIoMj7UJyu3oE4LNCb+I
PS6TUm2ZKBww0pLApcmkCShg98QY5dh4z9NzL0/xihgaZ1ln0CDkn9qdCYkTfA2/2lcwYkpaP7tz
+aZ6iBOFV11bZgRJxu9bsJ/IcwENkhlNuxfZ9FCSfwjIkkUsR1S3jxCKqYPRamS0UokjOaFm6wLh
W6M2BUAL7lvSE90G429/fN7gi3HQNn7nEf5AwmWUV3wtMlmVlNtDeGBWXwU2aVu2goOfIgRV18Ek
wNa0TVtZ5ojRtX6LjZUVm8kpU0vu9gWUk4S9v9PmvNdMIDn2YRi0yaiSnw9EX4JlcGQqiyT7EjwW
l2m6qs/QeP4dk/UFqrX8F18Au7PyTFNpjiglaalP+IZ6/FHriwVZYgbTN14o7F8wmd+GUqpD3R26
xqRPDvz5bCsHNUGnZeDGCpCqIXmhH1qDbj0xDrtdsBI3lxun1b/qvZkaylPRUxsXqCV1IIrfmOGF
stKDrNGjsRRYnEK/c5/nD+ceIsQnxpLk2IbBokyPLru0SHIzzE4YcVjww15KDBM6NhZYn81Cc+Q3
trPuAMXhk87VDOKrxQrurzd9hplrx0YSL86wGNbR12V87S+WaEUy7E6iFQSyHk3pUOZuz2kruTqi
3NfdCqCcpWvZSbESjhV8aCwGGzN21g7B8eYOxBK1k7SDbvhzJ75y259iZUbShk9GHyOobuwqNSMb
dJ9NUvOUQE0exbuMtUSnwHPb/KxxtNrd2BmVxhUURYL+vdty304Uc6oqfmP/ASx6ePRaW1MoIl2C
V2qLvczsdQc82dCaF5m1xBF4gtsyj0bqRhWS7PVrmMVOZtRKa2d8RFne2utdlEvuarsdL40pFiHi
t8l4Oh1QMgAwjlP5hqXdwXW5Ey77WnjGTXW3waqH0l809o1bggy6i4LgpOvQPCZR905mji6jgYOf
P5dVaNsO20/DPes/ay7EPNMgqBRj4d8LQiuFd0rVxmi12Dcza2r2YaHIGJNeTIrzmiRPCq5ZkD2i
/fTvCO5lCxGRBOnU2voFeqSnrWR6nQR7U3IpRT7dvg++2vZ4l5p4qbdio596/6PHizk+S58uZ54/
e2jPJt3DXeiOVI/5cmNxwzE2l0FyYHm9FKtJTcEosXylFBuWdvTu9Ky7I420e+h7N3HoEELJjnDy
q7z7h3kfNRfC9fww05tlZiE5vbcCFDgqqqpUbVWeWyf70BtnPPeZpF0iMb0d3zns4a+KfQpq0f9a
ZHiTGKpD2VLHkWJbZfabJrq8ZaoyrAP+nf0IHtDfVB2WL6ikjia8biug5WKHcGAOGyRj/v/vni/O
044apXhQPztoLVZ2R9MkOJyHSm1IHm16DolFiRnsRTMsXPAXdN+UjcmzW1WDDUebyjaUQJnJCLLl
EryL7B7jIu1FqczEWUGPyNKc3/tW5dRfXoNu69jdzp0clQezlyx78/qRBbzh4rERmy6iTFFyC1Z6
p+WC8KsOnNvAKF9G+F2LYNa5NrTnW/IWeR9PgysFN/KKAjlBcSLspm+CGK1ijMyovcNXYRQvSBZ0
X/pKJuRpS8HPIZrZZCLVTd9tUB71hh6vpiFq13MFboMObHR9A4nX3bOVHrb6hgHnfz6m/1R5Abna
C0JIoL+calUl15uFqaPXJmxKPz0VEFy3uYC/p846tOnv1qcT3pyDuQEcSeHdbQ8xHmAQHQVkmeYk
1OZ8eA3cEJ/2wCcR0pwrUDX50XKfYgFyG0z7ID83RM4y2evwMXATzEJviC9Sf+FZ2qWtCvTWsVwI
H95p9N2md2VB7BAtCTiNrXt0DuPMc7zymPFM4FkiJzEw+AVegoKYy2DUzadQbPSf/gkDueTuVJ7S
YOOLqcQjniLLgVwUWVyG9sWXSSKHjKVlaPO6p+WQrD9geKsKK6j/sWlMnTglvpGoLHQQU+TcyhB1
gHmXKJ5pp3e+IP7grhRZl3RzCmsyO7IvevypudW/hiO7B5menJrSZgal4tBYCl3DTOn/FRuj2mk7
ucFSlnEAFZFSCQO07pd0BC3hXmf4hLdTWP4i44Nqxi5vRJPf38OB/z2vjO0StXrS8e1ZnLsD17Xk
