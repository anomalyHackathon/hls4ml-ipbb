A3e8bBlYGURshXBbnEdU9hsJB8M0khNx/vlzVS8Zm+5YKITC3jFUGyYEdlk+Gjnurmc/kPaQzl1X
2rPSGpnodsmCb5l5LAl9XZLA2ewABMU9w4ocVkZ0tNMlQ28eJ1PMJIwaFqQaPGD5ZytZFGFIkAbJ
HFa0N73+sVPvmrwEMLv36a5FoGzE0gQLZ6bJW0vo8rJZSux6N6iZ3S7E0SZjwh8RqDzHxCDDlkQQ
bR4ZXABAQfzkKWxfYuK7aSXfj/BFNBV8j5U4MeDF0RVbGe5XeoWiK/8zUWWZGl+INTY0h2MytSSm
+XA4ofuqkG4DWvesg0ZPB98ufBfCazW3jDZ2alAYRSzpVZB2hAvyE/o2yG3GPASo/a4HN4LPSF8d
EHdkto3fac+kd3oG6lQr3Sm/9dZXjpfVPqyfqMNeIqCXfBKlrUKOVvUj3P3XuhZUgFBdKnw8atlR
YtmjtFflcaiaZoaF+YIHJvnNZClXMmTXN9ZqEjMz7bTGZLpa7UwNHD7uNFPGxCb19GcM19CqNz9n
EjP16TRSEjNPF3q7Zy2ZzRUaXO47ExAKG0fY6F6KOzxteGbgjA69jaTDxryHF5xK7mBTE161Z1lg
H1FAFvf1IhmCuO7+hLb41tmJoPdp0evRVLIeErBWxwScBXme7Q/UmnpCR0a5JyEqiVIPJW8U8sPd
7egoNapgsgkhVWuBDT2a6pzkEWeX/LISaIpTCm9bZY87bBMeleSMqmQawe7n0pkg/6hsAFaa7a6t
H0jinHsT0Tb1y1CLmruCa47f7WTe4ZYa2szYJ+iwPTYQzn+ndchOlMRfZjmGk4exNWKiHmvVxy6o
Wr4+ZbkyBZg4wVlCm63/r4uAYvLDBJVJqAxM+xaPpW4KJfbmoImeexL4K3bDhuiSGAWO8NS6+aN1
m5wxO7U+Woli/We3cxDIBl8K4QRD5luXC2CWaz8ldVKX+wmLTbOOB3MN0y7SuqL58r++80gbckdG
34e8abk58H1Ba+6kG5cS8SJGmZp+RuGb+JTIiKQeGdX0U1iWn6YYar8KEulg69FBcDYg6V7lAbLA
Wr7tvCgGsz9Q5gerVOCtuTA5/oiu7J679NyAxx+iiuUfEpzBrHGZZJNpLCKoC8825ctusxcbDnCd
G9pWPDay01jefEORDPuDLIAT+OQ3YyFGzH3jbxEmkO3sOsxrCxAYexXcqlyV8nXRdNBP8aEbbjCM
ZVpfKCKgklr4tYcqG1OS0H9IsnI/97unAHjoXUHXt028yz8G2zxwlzQUra1DWfcIELPpTsFrCwXg
//yU/bNDxWJw0e5cBE3v15u7otq+mZ68bnw5VIudpwwG9fKUoENOkaeZxvNy+JHZSPNlQ7UKSYDc
pA6Um2rCdHp/Uh8MEifQVMhAycUFKC4wY0mpqmWQIYJzJsUTuuAPOFDf5wZ3C3pblch3aAUaF/hK
TSgAZ6MLWK0s9ebL0oCVxEhOC024BpXZTO8N6Ya/wfYF+GzJoIRkEJZvjY7MkiuOUQbt4v/gFo3f
aAliP8jXxdQgx7pWU3t0m29izDDmLkBul/+efRM8zWp2LsNSTCML+Yb3YjBH1D9Z72Wtjzt7BBqe
MRb+hv8eL+SChz2vSCxX7Dw/fezqGH0GJtzNeTPE24pV/53JggMziPVxKCiG9t/qnp7q1ioEgeki
GbaQew+hwQ39SIY37TGLYod1vaUuZQAfm4TYD88vM+8EBKRG2DgAo2eLl7KydXKkDe77xJdbZMYK
PHEQ65RlEKw1+FgyKSzFzfs87BLy7xvO8RFFofdWAhkQIa3ExOJAdRqe4p9cxj9dYB9GOM9xh8Xi
z4B++1tEMRyyt8FNWKmsyp9071WDpg4x43N/yPkpG0XpPL62bPYHeFyqac7zk4ZnIGIfAVcJJfYS
PbyAagLQlnfWjPDeo4kwzD6KBe38/6vsCQz0edqjKhWeeehr7NZmDEpwwStyBO1Q1IpIFPtPvNlj
H5pPSFIAPEm/AiRLKk3C1ianahN2pSISIVie6DmGqYfUt5dzSb9dAcsZ660xfsbW3Vl48G1ct9xg
FEfqmSAfqeIfaBIqOpefXg6VfYWRPVp9Hs4HuXuzkE/r6XqoGTFZEcRgHgwbbafg4jRGmMhwz/Nc
aJeuFCoQaYGOZOewpxPGACxckMPcDhlyz7n1i0YXCoiNAAccqc884sq7B3FxeqlNXdnuQVfqolvl
LWT9VX6uL+4zSKCsud7YVTK6fP4hGrojCK6Pr4uX1O56fVAvfvdyH8IOx8MIjdi9RtDtn8Thu2md
aMjfs2BotlxaIOUPSr8sGIKt714+8e8WTuSqBBxIP9brfnZTtwDv9ogVuEOMEYZEFxiUTxAJS/wI
izhrkVi8poi+6LaTZXioDhHZGgBkarBXukwCYyXAh08mglhighVIQBwnHYvP+DaGQtnto1HXPi6M
qrVFXMD6te8tFgXjUTuJvWGUbl0Vg6uYo9M7//arMzgqsAy/DguDAFlUktSc6FmQ/3b109sgPalt
Dm9nMlmApWSplU2BJ/3+/fFSWigzMdHFPUBvfsx2RhJUxdk+qi/XCONBtgYeGPBeOJ0jVnF67KrR
pOxPY23yibtk5dOVrDzGimj4Gedwd1ByHKr/QFJDz44oTn1vEhG1Ty0Px4zW3OvlAbzhJIpR7GXp
fxGzHEWy03Ix7ev2yYDcnAY7wUti+OsRThLbB6epPf/rfrRcZ9M78ZBThNhpFhQP/d+nkK7+o4ll
dwtKks+I60Ys9j9Un5LsxdC3o4Q8jvkPHu71VkuMSj32D590cfnIIFG6RZZj+BqxiEdAopPcLkol
FXbtmvvkHBUwnOAnxpUBDTEom/Mt/or6jPqFaPCWwgwue8lNXyGhk80Rci+tkAlSM5etXefjVLB6
5/AfrCf32G3cKJqLvx42AZDvTBhf0RIDwOmkiftMhf5bLg7BoW9M2VgjGjdqcLUIfuTWZ6rNmZyd
FKudNyK1dO2TC8ysW6/EYL2WzLNy+BapxiVYxiJn7AeqPMKW73lo7Hajmk1NBIYJl4gMm0HkbOtZ
hqBK7kBrgDyHhrm7efCW79gLLA/lk/+AL93xv7RVzh00crKmLO/WJzVRu8uDF2kC/1/+ihqSAfOT
sDk+hv6qXqR7PXTPvZPctA6QZF9L0s0jaGOJDqF75R2i0MVRdm/NSedbys2wnkU1eYvP70UO9LNB
roRQlk5dNoLAvBIFXp+qsjYAE0QX4aVyaAq9C2ATJVr0/RoLak4PoBnWYE4zO410QwcinaDwSDwa
s5RnpYEr5JSOfh2f1ZlfnPYd842RXY74/qXFhmkSIDKoRfK8GB0AxxHxttc0TlHyDFrKAjcC6yr8
uy3DM1TlcpzgwucyqmGtCnM9uPGNPr9PuGv94Z/Zfx5kcn18RjRYsQZrCo7mGO6T9uC3Fz23abJu
oLmLIf0BCgvw9rR4kfdaH+Rme6qtyuuyVcwTPTvDNgGABxAr4vQc27Ps5Zft4+aSz1gByopsNAkq
dX9x2HnnmxlVrmae93ee4LTQfEIAr2BL8v9LpU5ZDi4XtpGArvyNkZthxdZq2KNkSb2KIvQnjNU/
sQwF0Dk1Djz+0mwK7XGhTc5lDTc8QwCIJ7SH3GCv5dfdTzaCwc7q3/0uDoJ1+/21tYxEXbnp9YdN
f24HaJvXr6ncyzMX/YnQEzPaXIHwR+giFDiT6H5JhyFHwRSNAce+SNG5EE/gBg1QinvwWDei/253
a0hjizkyHHt2JiUrimmcKMo+MTsOpfY8uj56pGTskrihPwgXGSBDjmhmUnCqxzZZ4pl6OKNxx0yy
cdUOfuh88LZsxpOalOtjd53xewFSN8L7wC7REDj7ArUVvsA9u0QQb/kiNDpwIZwe8cuO+KJyBepj
nEinFOH7phd3WVdnTu4tcF2rviS8ym4OpqDITyBM5hVrAj3v1cAIa4SbOY277B7QxPlA55nvjgy/
aBvmV7AS6+JKtaMJNaiuEu999rsIRjQ4YYXj2XfLrUNjfAG7qfiLgSu5dR6+uCx/DGUtSHIyJiaT
Mil6/6qo7L3nNnceYs5+0Qsla8ngDIFz+Xuo//T7bxZK6pJneQOtogoI5Vv3y2lxpeh3OQj3z91q
66I4fbn4oavQZmDvhlO1YSmLShPM2Unb6WUEZ4ttwske3hDnb+m8/njw60SdLZZZlr7/c4O3e6jP
IAN/MSu/TK7PVTGciitq1aIPKb13UzpC8VR0K47X4LaEiktYjoWi/YGsYpFg8ke034y9oWoirsI9
g8oJCFyn61dwBHAP4Ry3aB74eizfheDNprqhUVOa/iOsVZ9fM67tEe7o/WKCQ4kgbZQL+MQiNMyE
oZ22DKb6LegNf8MfKjejBoPwfOd3jPU1PeE58yChvCtNfMz0ok4X6VfQfAxfTeLBK4Ezw6Yl48zj
fyDw/sjzBohdSctOxxpmT9dbsvlMA9sUjOdA3iHu2hxyZ00FU9FEqdsA2X4azttrcJvsgfy7DRQ9
amrRxan8fFxMUbHxsV8vxcGr+ZhaftWicge9/D3IYdOLsEXd1BrDQPiIm4aXFzxxzk/YA9dZ7/Ie
0ncZXMjgoqwgrpHIxmWMw/f1H5p4YQTaYO0Hm86+CgvfDjoqcVLV2iOLsIco15QN1y7bGl3UYH72
dSXlqktf7To3TlK93IHpvR4voLwreoQ9eZMIuhNTS4uSJ7MZCHohKG4u8gHjV+wLSyAu31wfAazW
qCKeFcJQdWdbr8X2Lq//LBtifmSmklY3cxF6V5zB138hATyl/flqqFXNRm+bByt3vM+iauyeFRqT
1G0QaduB8IlcSe5l8Q5gLlnkLvMJi5xWA4iFacX6E7Kze/Ywx52R2jjDO5G2++Xauaq/P19FraD3
5trnBNDRIwNcdbwESvmXZpaZKlMMuOTBw69w8tZYGRLmvfGkk4hTYeQFPqlX54zUt+st8SoeNWJS
v7p6Ta+RAgIA6bzo8v9RcFxMb0KKCE1x3PfpxPg9nPttstXE2UKFPgl9+axS75iRnxiJgiR6bWsl
r391REscggnjj8X/rIzR54ePtT82gdbujANJjanstet2ftZi11jv09hMImVvs9VS7e4Kf+yvjv7c
2X/PQaPj0WAIprdASP5sJE9cn2c4dtAchG6Ylp2GfAvVcrR9bE/FUo7tZLyZHlUmi7SOrVJqDD3T
vqpNNghfjZioqONyOzm0nBR8mR3zr4XmCF05E3C7ts9LNxArHAuUUsmPt2c7l8uDrP/N3kO1ppca
1Rp3r8mRmubbvos/ouk8ZiYN3IbXmY4ijl/v5tvWKLkSq5VOmv6maJMDUBS25pHjt0hPWLK/4ieZ
M4h8FTbNQ32GChgCJW7UyAZnzKMTsVWb1K/a/QlaRHkSP8J9zYxaXM9JtURd+qMlN9xqa7x/li5n
YFaLRyzVratSKba4Cg97tU3JVXrGHgukcGhmitG8CTQ1u1g4J9oH65dOaV/caf48XIkjZpWMWp7u
tAkIh3fCKcCohgGqYYEA4I58mDrM9u6C00oCRJaGvfclYxSl5uvRV8IDAVbSRWhATI+WV2I6fdXg
51NN1dLP5F3qzLecNyPXWREnmKuBPbg4XAzc8EGKEU8jWXE/TdkYC5yclaJAKkLP8fwkAqqXncmW
6hwhcTZ6nzJj+04oPpDxR4YOWiIkGbZCXhaWzdcj7cU8ntCX++2rKqWGhowqYFSC+z3tnPpAL/ob
oJ0psGIq5tXWv0hnacstH9lwxN+pyksX08fGuxu+d+qMubviq4jRniPszqCneZO9v5Y1WvYHM+AN
yMeJwOvnaAecvb4BPj+1CrTG32IBaJVyMrhSoQvETwZFM3Fn2yomcU0hidGtsSdnYdZWwitPNEBB
IB9wlSnYblqtyay4MiVlYl7Micv9IyLXG4TRhsIoRqFKBwWs8EzNoU22qT5YbVgowwELqcFrJGC9
hwL84Yj/J1jtPl6wN77bQO5RH8PoyuDZqIKkeSSu8iH1YoQ6QCgU/s+8jHyDOc3f7YqEUzPNFObx
Rb8X9aZD2xh9sXfdsS5tIdYyia21SYtQ1KBhtAbN3yU9iNLUjhar6UqZXvbn8mbP6sIxwjF4lvhz
5cmrEEjcMvdY7QQqgWHu8IeNiwr0SBZ9scA3XYqenVv3x6YKX+AvJqwmdTAtXDgvBcoB6oRnpbV5
pfGgy1+qrBmrOQUw95dnm1ZoLYE/h+OrY0+nQS2Hijbn/J23azy7+/fHSTx/HJAD6s6nWIAfm4cv
UC94Ds8A+ZFvAH0lQfcd5zSd0/Tkm0teb7ZrwmifiiUJYThiYNmMpZ68W3eFZOBXO8fL0Lj4PAsA
s5uUmT83IA9xAkVCycyiA27GRANr1xeJ85bmGkOi4l3uQ7xlQIyorQD4no3OF6ybMJhCrlmqb/sY
86jDhbsgvuDXHrjU/CA+dIJ38oQZZEwKZ8cLw7rPXnyoDIORJON0wgd4f+vQEX71FxFRUlbUfI9q
0V6Iw7luil2GkCOhOBFgx894cTqKHtLy2iNteJjWe/iBaXq4VOqNlZ+zpUYbzlzOQN4AasAabEXh
sxQbcAIOYZFYFWNp+amuns8puJo/ac9Shx4USXBChG4tTlw78VDv8YjQPT0jPjDM8wESJN0hue9j
zQX60EXtUe5OJOQlLg0tl0N3WMpnB8Safum2sm2EeqcfT7YmrpHqWxJIb9GkPVx1VlRVS05tMfOA
apP6mQjRLaN+hahJokt/CaGJYASpGL9Dx7M+IH5XyfgeB+RHM2gwEhBA4ueQo7yW4fkaN0enJMSV
kwLXy/q5pibpYTiJYclqi4pW6vck2kIXCLqC5AxMWZylaFMM07fph4EyOTpqu93pX/hq2vWmf9Ig
5rjoFRAVFB9Tu8hYUAhttCE/ul7NEdyuHfjQ/mMD0V84wrsAmiORjDypuJ6krLY1ixDv18rdovjn
nxA+Tp3NeTI4Ub0BYQjzUw/psHc+5HUpGslJ5AIUGaIbZDwgZfGLOqJswBYRUT8V7pEZJ7TVGvYN
GUgGXXQMxaiKPw63wzyRYmlWvMLAwx9CB67qt/w/5DsdKpcFZtMjWfo8nJkUcz1jQ6jfzYpbaaOD
cw5J7aDco7fBlznNh2Ta0gSeyGx0zxo52gRb0mAigne3oAj398N3W5Np/UjTL429dGgL2CM+DkPR
ZCJi7TrR+BxLLchoJdK6aewqazVSpzD0MqDmegBssy9Djy/ppoMO6bAMlUwEivTpDv9VSgucxr27
6WBaWyJvhLrpo6yymYH2qq++xgQfcM1aMG31jKgfoE8lwondJV45FrpYk3EqjOYIKsTtMQkZaG53
2akfvCdgVhjqC4XO5MH5hAmjsbfHIQSpKD2Qyl5/3om/H+NJBHqXM4Sogg+JYuQFCIekfDHT6hJN
uyPcKIYQWMbnZuKfYEhth/9OHbpKV/FqFG/Af+mkCCGCdnp00RrChQwfhMLm59vlUBOWYK5FPaVt
zn/5LRMlEYDlAX3IriO+dnM58ccQnfEjobML+7Ad7HLZqxk4SRWOfPPE2N4XDT3jCRkDYaa2HfTR
NhXLdWeBkv1sfUJfNI4wk7bTTzXzIxlKVxxLdbuqWpx/xx8uD3MfnXjmalo+/j2P9oUzO1xbkiGQ
YzPrFKnof5ZqVg+7t5cc1R6LxViaCvRaZ1eZ9gsN0ZiQRH9jgLBAq0lFtveNxgx3RQ1zLtFJ/zto
kteWLb07vVdwj098gToETwCyIm6+y1dsyJaxa44XT4kGoAHEv06dL24V8/bQNFvEDjBSM5jVXqPh
nD2aIGtLrq5/QdxYDT1BcKUqBZeaE+EYI2tbWOcFgC+9LHiUFJuKIAn7JoR42r5eqQU+lGWDwGVi
uJZfognJNQeHxKPRXLE+hXAODTOVZimVsWBa+weMYuZh7vy0gsNRcFTXfCvW8g/SinonqsG+Trtc
CEyzj4abJEpq/qyH4t3o+VOFtcNxgjGsi+4o+0vgE+Qv3u3jf8jCGLm/6CWgmF+vMFv2Yt3Jv7eX
sRCFnBZkAnkiNxx06lQtlcbmQ8XTbvP3kiT5351/yWQAs3TTI3MnWPRGZTdrV+UgPcr8bIMc9QA8
umDh5lUG0i4pOZ0kwOBcMvciiNN4PcqQ7qkOPglmg8z8gCziP2UGMuF14fl5PsbFbWd8WnSrJdk6
HaCrUSfOKcmX58pgGP88kLz/BW0fHvhSVeMbjC/hKWOvjks0luk9fHDipwZlMLHlrmqrDsDvB/FA
1y3jUlE4GgFZ/MP/UJTRtneksuqCo2i0AWgYnf1u2xizN26RwoI2dzJQ6ye73rcjZOVsQrt5u3Ga
a56njgSn3QJop03qRlgH6wX9boIim5iXHaXpMPmWSQBbUmwzUWMr/e+/ZR6ey4a52UHx4x1WlF7s
6yCRFc2gw6RGybP9zphlnj56L7SEOxrovR2BXxPdIIWbTLuDE+WK5/52xZxO0lH6BgLRKhJXy5w/
IldIYPzl94Lrow3ZyWFZDa6fpvtLtMEzE22ILPsvWYMo3yEDOupTSOxKY1Bdb3FXFthADFsoTFDk
jt/CqwZPdyDccFF9taJMVrsri1yFUhEu6VW6nppJ7QMbIxcPP5GJQnsWwZy5hbB2vzJKV0ara56L
3WEjVHLcy8kT52bVmggxprR8EzcKYKxa0nvY/Swcr428cpOW4RuoevkNjX5YcnZEVJBD8Qijne17
cQICpreDHPJJGoRLZqjSAJBKYEyMoK5wj8AsQFOce+LvzU+Xxe+aj4H3DVcOZ+nqyWnpYbPwfyMF
lYGf/Q61FxDkn49CzXQ4Y3eCVOo9c4y1NQwf5rkuplInnld4EE4Ebgko05+4zazyN3LOf7NWsuNd
f3vQ/+6vPzW2d8lNtqZIgGtlB0Xk2oc0C3fMPtcsBBha1rDjkeSEefvKVcRuCHpEXQJZr7WADtBQ
dk6/hoD105hZyf/ukCZnd1f50TCh5XKCFqwnSjNm4imjmEKJe3x45TXaIYpw6uSX/08OumnlnGaN
lQ1FXilxHOsv6aw0dXFLs+qYfD88gkHhbJ1poCVZhMzY/gVvpUEZoFZJ1G4ilT/caIyGOec9EcD2
JWgd1XgJ+MpvqGsTBhzTfRVijOFwG1orpmyH8tcBYD9EZGeuWZpELgKw6vXj3wvCtip6GTLaK+SC
4hk40raqIRcWr1f7/blgKhz69weLMYJviYT+rVJ18L2Cqh7L4wxHGpkklFRgEVhC6d52IxG3G6ZL
xGO6ul8xH4/m2QDcj/rva1Izo/T7H9tBOACKHGTPawcyhMnvR3ra/IT5DRG0tI1bBSENR7b6EjYH
cE3YLG3wOLMjFsMa5BxvTUY8V5TX6088XlijGtTaC6lembLVEWQv0evEoAM20a02+AUW6nL6CJbW
eX7DKb8+v6P45ZjH41c+G6ToEfpQMxXikAJ9PSWm6tltQL3H02uvaxfiQnxs4QPfYknPm3bDUHzu
OFJHDTV7H0y3QmuBiErmPpDYFjez5SXIBcDD3HuGQfEWW7HU2HR9kTLirZVO+W4imxb7xNhMjlMB
BHEd4PUfw7K54SINfU97xD6NB8LP3ll/nXcEDgMl0H9F4VshUGFJHzscA9avsBdzTdTGmfASCOTN
o7e8l4pAdFhxNZ0AED8iuHJZ81cdnBIbWNPnYSWzoyyvGiDZAhvse/NsVk0V2B4FAlQFhG+8r8RQ
GG17fQcDKqpuNrBZUoyD/u6aC2J1rgE9TfrMgR/qAEY+JhCcXvoKsu9hMwGzMeajgd/582q76wlD
l4qL2DvOjr6tObIepuymLPtAX2eYgdO7onIzSMt7QcbfEv2Ts36EvEzcyene3j3fK/LrZD9wm5BU
gRCofdkkcdOsyRcLLwt5C4rme5t1U1LUKM90YTorpT+5ptCl/e4wTpDwoFklepmrRzHZpnNbDvAr
bubny17jTYiTQvSpT+TXsY3oxVMnPq5pwMwah69vFrfFHfjliFQXR/Aom/WpcSVN77xv0UxxeFfy
PAMHopuFvDbRwE+YPaT/RsE1uDQ5bmXRN299jjXEm/pzpupbfMi+s6q/8XQNRNM2xXPlv5F/k3mn
53TOgO5+ELXL1if11i0HVlI+6RnZUjJO7PTushS4uSOyDa6676NICIlKJvpvmAmDydNY2CNRYznk
bABxC+Pc1zh0J3vdIVY8CEBrk6Hdsu0l9bc5MEVKU8UxoIT8nog8zxKSr1p49OdUCy86KYR5eSO/
gq4z2WkIvw3b9GD+6+kvuowILZFd+0V4TmdndlhBY+oWz5TC+fRQZBF1Y1zTTpAYSgCJFiquh1oP
l1pEJjgMvS3SCy7SZmrTD4eLJrYCQI84EQd6DdfIqmTwFdPJA1fH+U6Y0BQjaqq2VtvVO2JvXyG1
CoSaiOlxW6sO81+1sEnNQabrMysbpDbU3ilrV9v9IyyFsLtyDx70CJ0z5DiYyvKVzAAn+xfyYMbv
Igppfvg4o7lm75DDCIQNkksxOdKH9Ni6p1W0th8v2f2mWm2yLhG3mfLog409ZKoiyRfkAeJdqrQn
OPniO81+gS7goxKTnSstqKyTUtlopZZFMrt0Ce8WsRp/H9a2glr3APoHxhA5S2w1fWl4ne7KgucP
KRtkjyp9WzpLnIivIwrqDI42eFBIdVa7ijQdyJjbNN+8CMa5InfrIxu8Jc+geSa9qEMhqfMTfhlc
qHLuJxnKVPgxh1yt5yakzhJjRED06YJzKbHSmCGtNo5byTbWT7v9nl5Gps/4MyerHL+GZR0lWRdz
8Gp9Ta19WboOebtqOVdnduuOMnrBqLuRP8WGUERcPLIOSixlVMybpcB/yJqt2Mai1EopK4lqa+HV
iI+5qTr6PHwnQmYJZbAyHXeADd3xNGB0hs1Ak3Qnjw037BKXVG8IBEfIIAGT2X6dv+LfspGBMqZ2
k/fZaLAvuBiKT+HUi/cXfrUgzUrbi0UOJUbpZomyb6jKGaFlKwawzRNpWaNXzgliZz8q/59v0NtX
sSwHtgcVKgB9DN2dgUKy2UyxBKTPzo1g8b7ZVmMxUVOFf3GWawSx5yM+FPpInVrHUt2tuWOZd3C+
ucLr7Xou2w3uO22VdnOqaa9olpQdX6dlJP0khE3ETs2o6WypsEFNXpaRRexeyqlGnVaKx905Yipo
40OefjF0QGbWFOFFOBhpV4lt9hRbPHWtT1HhWKY2LHaSjL4o0SShBSXTAN5yj8TQfUwRlBjrbEad
hDW1EY8r3PCvba050Qzd4NVjyfo575Aj7F1gpkEH9dBpe18aQhpB9D97CM6LehWZqODPNzWzBzKZ
QlFgURbIOCzD0OJ4YQME7JBGnkCVC6Im2zP+FPELiOtbqEHX+VH85nTjhH5+YVCO5OQkjmB0TEqW
kZHk4m800kdFCChXA/aE2RHJ54juPNnESCnpPBk1RqPYa11hK6fJbPTUIaqFBGKw4nPBNV784iVL
U1nKEHZfDcrIVf/UMACHXnjeR3mUsLIqeTU58Kjv2MSKPdQE7t/l9XRZY6QE0gEPo1kstIAYsPD0
EiKpff6fXrKKR+i8v750keEdJUUmZsqFSEIeX7cOkSzQYUsirfMzNikN8NrO9H3vjoA8yqXhUHHF
1Qu3c6OqVjVWr/509HAPXEIJkd/8l5D/v5bE9zcDx4rnl8OOzAJNROEAAKOwb/71gmKFvxorkPAI
RjwNEaIFNqRGrjUva5u5ALN+Y0fxbLTyr/FZdqso9b1fzPOCVEg83tq4FrKD9yUMSmUmI37i9qVp
R+29ziOLtITg3lJ4o7/8pDOgH2wBxEph3/D4lBoz0FquPnCwfZ0YUcEsbNTytHEtCOmlwe1p28DV
1th7C1NS/rSuvyUxNGn/02vurYJUV8rwHFvKn4HFCJ4ZVssHPB/RJXVb30Ec6mGQWMvgckUeETq9
hgSb2TzUKzz6SRE0gHFLaWk7JJwwKKMW3Kmr+Br6mdZj7/H9CRwfax2nM73KDFwVtkK4oRdHVDuP
O5LjzTzjpYSpdOLTO7r5yv5ockYQpj4L7jlBdPow3jtb8BSL/mh4ZvR2DafpLNV2Uf975fdC0xYD
jXOmiLORypFglRkKXxuWMnNDNaYg6R3B8NT0RGmFhuUfo21qcWnaHrKsKDJaV3p3/cNfEirn9YEF
MAWz2nGtdMLk3bnne+TKzsZxCEOBmRNHR9gSPaXJJhMMw0Q1M4mIzN6u7ywfs9P6hJa1uSr/3rYF
le3mXnf50t3oJDL0kCybVWAi+zf9sc38Vaku/7nbfzOvoGEle/JxKUKHSkCJkQ6X5g5lKh/4kAgu
++utE5Qb3L1OHF4Zkb4etAZsXeUUnq+7ghdGt6fwKeVMOc3ETAvm02m4BbBwAjiSUufX8ghm58Uj
8rz8Ipo+oCDacyXY7NzU+MtCDgQFgBzVT0vrn3KvzomEQHFJgpk5VxhOZqlV97FrfJtV6rAxiOnd
SMbtdQyoBRBsMSbLsWMb8kD6GKy6s2C/Up9ZeMwY5hxmo0jioQip9SyErJ5MwBWYxwEhvWUNti8U
LDJF3yckiL0kfpPZHAjdyV7QlGvpOYb2C6FecXmz4ExsIvyrej8FjVlgFzlc33bqXW6WQp607duP
habFEy8m7d7LVXTJkc76TVpEV/Anf7M9aCQAWabsZLZtwqpgDupDL8yIZ2GwNgaFZhG61NQLqDZS
NtZoyiRuyZz2Q5qm/ak5CTfky4TDSxd11zjxY+wtEUBeZxtcIb6V8Xjn8iqUOQ1ZYNxxDiv1i2h0
Q1xi4FXvLbknO6Kine8wFe8Nrst6AtGwXhOArH0eduIDo5LLdLiKmh8koxlaBgjxyIu8fe1K0jOv
dsJWTveDbHo/METx9/x19eHQAk+njo0aXxCDd8wn1DlTUiXdUaiaPDpOEDpMNgWW4ViTOL7yGpnr
JUr2l3MSexmOFfPOENuuEZNCwTil98qIimWfQunTjXaNPH7YXA7daXvHqddvdw/zO2vFUpdh4uAa
A4vnDEDlm/5tW6S6lZdYRDYakDdwyFWpCrvsmWctw8JOsZhOVrsVOqPu33362yBb9rnead2tdPfL
sx3WxcOpiF69qWSzP5oFCQBWOAp3s9W2QzTQFXMkQykBS9MJSeziw3Tol1Lv5WF6ekjpJM7GtLEZ
2qT1q5mUIqb9u9bc0R4PeT3Mu0v7YT/hNkH4lUGZXxY1RnBIVsxt4KIw1oetgjuuKX4DOVp1d6RO
3+hLCCyHT8sH/0H1ptO/4pJRT0hedqKgAAlhKib344K38ZTjeIsXsszBBasKwxbEGUx1hri4X0XM
O2iawB8kyUYCkNrwGUfF3sjOHY2FfgPdMZBLBsbqIQy7/5eFt9K02nyg+2C4Zp26ItGZmJ+SRHd0
sUw6F36cEO5sTaRvdA6A2dp8bncaGiThNp1RB7L9MA3opE68w5mhbzAMC4ydv4umbN5DJHkkVmdT
4s2yb+BNR9wzvY0OgaRlJK8ZntzYdcXXnGQjbsQ/L2kVgWXAga85KLj852SaF4N0v4fc7Ensd9oI
4sbk3Z9DF6hiQfAIVSmBYvf7foBh0U1Di7Nix/2M8qWqdnBeinsRKxk9qv0XyBOtuOPL1lrLx0V6
r3ZFMarT9Jyd0AkgldyWwTW/3lDWlrmP3Pz7G0DZyOtS/pDPKo0TTJThpyFmY8HDaqvhi1mjuyYN
WNhDuFxPQh9ebgrXQTQBwYL1e7/Y2SRxxoH+AhowI23PEanh9CVfXw6Fn+P5K2kNyJ/KeeyNZtFw
vvmY8+wGPkL4KerAO7ePJGkM7aAIAWUKIV825+64ocsvSpz6kJu70VcT6R4uqDrQ6N5jZRISBinw
2EBXW8ue3aGYo4x/u47SpaDhMwd9zPizMQCNN7g3dS14yL0DfmG3NPVtBF3qinBWYOQ/X61EXu4Y
ugAHsxK7cH4z9xS5eLohXDhG6N57RlB1m+U0+n9Nqz0Gvl9rnpht2oStjSXWgXzNGPaAZDrQTZwn
kV05OX0MQkzJGoeKSbNQ/+/1u228KUGEwlBlRqux74Qa9s21E1oFE4oELsbTrq7jJn7qDaP/398D
5Kzkw5BQ85/h68sY84I69mxeWV7uIM2SPbBkwpog/RHqdRmfp1f48YWWnNiEdWpKkmGePmP5QDII
/O+5c0A9OEuFjMOIx9j9rI1MRccMMiL75W6DSThaNkSJGPV9/Scmi0wV9XFhyyeZXYVKCJU21Twn
u1m6Bf0rc518HRbCGQrTUnrc1Qvjvtcn5qpQYygRJ2BQVE851qp68DwmEkyu8w+NYuxp4Mglfv2r
+tYep4teugqhejA9sRWkne4KimGvBrVtw2uJ2onlcgpc6J34diiloEZs8PtaABqlRketAiEIoeI5
//bXZ9qwnhPVplKqtPsTsfB+wIdRVQ4XU3UthC+iOzNQxuxd9v1BNgtgSh6c3tNBUJ8S7IhEiOZO
4bJXmsV1b/lySSOmK+VULRODBSDQZSLMyKPnwjfvPH0HM0UnrzT3nwadfhd5LY0QZBVExHLvMwxO
FcJBtReArl/1NYxjUv5Mi+/XzyTG0kRCHJMRgrShG3A0S8TA1rC2JVSAuTjqYBi4l6yzNVG71AnY
l+BBx264ikOxGd/WVXq3+lJm4pdLpUIuxTfNZ+MRyfcCsvCAxLGifdjzTb3S7ovBkJY4J19E3r5a
cK9sNCkvuZgM1W8tGkHVygHplNkpBrd2+JtgoVIbnpUsPfdMnBwYUvk+xSe4c5usTyKrlteVqFlL
woebUkUMRNiA4CQPrIyOvtfWVwZHJzmyVyOJPR6RTFnxKJqEIOQpqPzrACiPeqUP31HC95sBqv83
li3r8T9UHSPxCk2PeDKjLx9nSF/inMfY7aHlueoRanSsKxMc6fGe7AQ4O3ntFhDMgwA3CYYNeLNE
nX5DcwxEkgKBRhSYFeevWNG71MAxY7vzCcx13Qj36v4rt4Qpz1fRs8P9li00Ilec8hcwtMFl81wQ
3B+2h/clX3pd6wiXgaK7Y0TOugolfZKIYBtimNbBzfD98UK8vhnh96yVG3rte2J/v9V3Vk/vRXS9
UVRetKEGLRCwOBE8aNGLDS3aghOm/WG+WugTTCl0+qZP9qm2GrtW17glzj5Vr8ytBHNCThbNkHM2
Hdwa+BYPJzFBv5xLSHjHiAJKauKAw5nddwb85ERuNwn90lceA7JSTmzDXEo5hX/EWY+Zh4+NFx2V
XrHj+fH97aINZL3rrMxUJ6McQvvHxlAUiXj9pT9wqQYcabKLCuPqsprijrpfoW0JaBtzFwlI8A5b
FYEF6qDLhNSYl/obnfmIO9W7RB9KXuoGA+/q5swyU6OSfDktWWNoxiqQRFVuFfEW2H61VJYr5aRM
ejo0NyyOYb/B5tqzsBZZYe61zoR2WfuJ7qafBX9J6CBsB2yOeqHoJM4ESx0toeRwfzz6PY+iW4RB
0TeMmPyjOeFu3kH2625BgWLKhvueIHdhz/C17yz03joFP8oZDCg8LUNjA+HoXEe4vrwqVFZKx0Co
/O/fccETaJOO81PmWv5ZvL7maB2uqaVhTz9Mn24Q9CbEUHe1nS9BdWy+Rwz2enPX4/4prpG6ZKmG
/6+6TTnhLgb8CrbZUD0+9x7yFSyYxvdzqSOT5qWZ/hkU0fMTsTULxtVj2tgRZxinDKK2S5ueHlH0
oSgxUooZ1UAvi8yMW/d6MJOL4LG1AECHzqqhG8Jr4ybbNWSEv3QaieiTDRlbqp7GvrNEVIm+I84v
PutVVtXPmBmqGMj3IjfhdqvtoljPe0BqwYW8LGMvpwNwhKliYPSjYAMkqs397allQrwGsWRXvaVm
zr22U+9zGaIWzj+n2fpgKFhrDewkkijfU4Xbxd8svssuMf8Cuyl1dhsdI4meCZgWacxSFpHFe0dj
1X6x952pKoK2McZOfOXQKfa0BSTq1ZbdC5N43lFger+MN2jMPXuYizcgnX//N3UZb1qYz0En7MA9
3OyTlh/iX+lQmUSsoMKl8eCQFm3uyxieKFtyzIAiPp5chl+H9CqQzxzg4O8hHVhKqquB/TOBHC/F
qJhPsfJAtQLcf/clcEhfG3tl3WvEBEq5OzLIDbZA+ZTuoLfzVxawez8cS8HpqdFNQav7ErkmQ+Qu
AM7qWsKoXgq1kkKlOSfu1zaLeETzc3hvn3qWAMOz+MoxGrQrdDHtY67o47Ogzm5jNAr3waGmAZPH
y28/GeM4YVJTfXr2bjsa9V2r+Cas7n79f+M/UxhBw+r4cizeTLTSy0DtD9PF0JwNNVne4MDR9a/N
7PNDsvM92cQcAv88shJ9bebfCcZtQLn7uKPVR0qGvnpW/YnHlbKKJf8RLAxvp3fMoHZGTK5dOqNO
p3rt2sNT5pxWyJntSKdoSVUhyabbtRGpGsfsLAjlbQ4fDenm/1L5DT9ImoKxW5lFdGRSajCfzkLx
ZJHHGyU07y8aTseMrYA6oYRqQ1pNM7Egti5uuuCC/B6/YglRE7tDKxcOvb2N5FA04vdEVflYkSqM
BLXuApNjRv9ifdY7bhS9qvJj7whP614ELmfYldixd7sDsuOZOxFZZQ+FDdnHqIuSFYpOK5y0/IJo
DqRfaI3PByggOAjVxjKUxldC90cAtiDmEoB+61ug9HeJWyuEm2fny1c6jEpamxqsmMbp2vOSkL0I
/Tx1ZLh+v0FiM4obhY0v9rGsTOhwE5Gdz03mD0g9/3+ezL9JdpI4B2w2DM6vOvWvyfntxM3/sfG1
8Vye3jdYmmZuTGnaxlyzML23xI74W4AgZ5zYzW9lASPOZ6uh/CkD1YMx/6+P+zQHugJK8l+IbsUt
uYtJ5hDLisfY5V9hx4x0gC+/9TN/i7Fyx8kcvxyqtTPgqX3mmZ1lXlO5IUP23Ck83pEGom35EgFu
DOCLkAg7RVoNKxCiey9pEWkZNZcVLJ5WU+jWBHWCM+Jvfwu9WGNzEtVu91vxAHMhyUZ2QSGFvjYk
rkaa3vkOZN/TOevVIFUqWsM8frMIuy+QYNXJGnL2QIqhfasVr1yJN6ghD8JVmy8xVfupr06PLwHh
2JddyiKdIxqdAeKLoyOwBv6AISXtSCHXwO28o8YBQkPd1hpMj1zthOz0B2dLTkD+Kbs7UIhAGkEv
7yrP39pgwGUYFo3FfNU2smBgm1QgR+Hm56JxbBnvOKk+ZmwqIjh71eWmWKqSvHalGX2CtqMd33wz
ZSX+ApRO0FrqAGwOeLpIm7KxLIbJfCsA3t9nc+nBA4QejmemklFdmT4OmWRhE5PZoaF19oP5Uclm
RHOeKPzCmqR0Cp3ZuSZ2mJ0s65Os9M3YkNhiX8Xc5zYXif1fykcLjO4JlAE7J7Gk7+OICEhdKsWM
vrVETLrCLMeizl9aWO3PMHWmsfowbEr/8JV5PweASRQdwa6cCpFtOq5AwX/GpK9mTy1lzN7jRKgd
mq641p/hewweQWiTzkmQJGMn2OvFsyMYOYi5wOVFtTUAidQ0LVy1nhKS5GpfjivzUcURbNRrxzk8
fdFCzCWZbOP95uajkbupKudZRwvao/qspCgZ8MAT1zkGvrfOcfI+OD6r9JcUcfmlGMQoypXMSNnt
xV9J741Ql8wqQSQUy7sY/km0CbFNmgmnQc7jevJr6bNl9TU3Nuz6NVAkDmfHA0r4cRMP5e0I9VBR
I9pOlrpU2vwMBUAIeBkjygSE/L5GNIOwGpX91cbJjODMreQfIdfh1o5idFZ0CJxXBimna9AGniN8
hUU4iIrIUjZutvTvt7PZ2NwzxZWF60BR2zs7l/w84t1EEWvgBspZaywTmt/n/vWgVWjttbTa3K2j
kYQMbSIFdDcdYLoDvXehQXefqBZBa6Zo4fA7qtLIIu60otzWTkwfBHDdG7jJGlykwM+6cUZQ1X1E
Z/nHfe2TDU+e8i8wpGK4bBblsvJfInR4/aFTpl9HRnex5zpc1JJ/g6TpwsNUHVuM+lhYg5kKl69y
ZsGaItvFJPIV58D/Aveoj+D4MNzk4VWzlx6fjuKWYvBwgKt8HYMJSzVUr/t4tHl0TtSz/p6S7v8q
f0AsmfjSOX/VzpFji6p0lfy93FYWVpe91Yo7KNMx3LRtw/dCZlcocq4Fe+91aIecUxS4x1Vtli/3
xokDa24ffnmXwuUJ5Md7E5AjfPxCsjgdlobAP8XFjVeiA6SnP+LLKPWuitT6+tR/I7IKFrRlJv+D
vG7B8wyZ5v4G5s6/h+u8cbCrg6Azel3qvdCbCbLZ7OGlQTVuR4ZQsJgC+L8QspwRTtJUiNV2e/wQ
2UvLMgGIbOAsCaAdlt/5ra4O/XqGiU5lqTKmsTY5j6gP2cMbn3ccYdwKv62cOJIjD6hjPzYk9tTk
ti25bq7IH8u85raCIzV28pCyxKcsdnWRPHhOWYLrFLJpYjvC+Id7nav2VdzxYqUe23aVMEm4Btfu
7vEoxmbYTlKnmg4QRFfVmxHHfb6tq+PAT5VAZRZCHng8dE/RHpdFWX4rADBSN0ZAabrcu+HxGUed
RFgD9WSrbGmMTOMmGxHA8XB8YA1c/wf2vJwnsBXRxpaj3DWNrnZ2/hxjKR86zed4V/67Yj9Qtmcb
awBieLrB+tIoI+5J2mgz7yp5VWphuliplAn9LD4mC161YYoA3cExHKsKujRu82PHE0j8ASvRq/WP
eUD05nmNbjaG0IVEsZT9XU4PuUmfP/GpqC7wtJOXqw71SgSJYsG8ucQv75LQqD4fUIJ9ZyfBgJye
gC5TlncvJnwdVBVXdH7zE7n93WmMwJw+Q9sd200p/CCdOKotdXZYilf6QcpBZ5F6hXiUBVAbf7Nq
PgZg79ejdLmCEVnnXQAAoVvpDbbiBDlRdiC4R4gi4MXr9YNMAAsaHc8EqlrvzEFLdlHpAQ0UxKMH
WLbMVYw83VaRJR/Y5LP/cFjLo3JDxmBNzWmZrxAJz2YoAObfLu1bH/dF+ecaDlSX+Touq+KVGxJw
Q4ca4qDnPYFvc7Ne2vz9wfDAlnKa20Sy9ro/XZoUg7h5yw3DfuHtE9FrSSUr5bZfH18AD2Uostql
hnmZ32T071Mv1g/5KPY7cBvOtzXiooTCpoOqZTcLJGZWGzvQF9ub4u2t17xvsnWnZ/aeNnyTau/T
8yJjCyV/dGOdn1Z5mEV6ocbh2pPOgfcNy3YBF6FASwiFRBrh7Qan8adxqYy3mnv9xwMVfVCK/1jE
NDYKv3tOgnmGUca4FqEVCwnXRCdle4Rv8gYVr4S0V4l2ShLx9+PsMyyYNuYV/DN/IXvrXU3bDInX
i3T68YdxVwyrnGZdaYSIV1g09hm1TVSna/lM8f+g3F02dlaQuG/7e2w0+MoxGDTIB/x4iHCIaewm
oSr/UnLISWK4dsyxire1s0vTdrUgye9yKZXPpJo2NzhUmBPBtrG4TISXqp1udrqP253BVW6PDJ8K
37/+J0jrqp5ZHXn+KXC1kLLK3eSVOHTpjjJ52IbGH7cjhbqodIRYyoJWRL5dNmtL4MewzDozXgAC
pzkuwps9ELmiRSHmSNDURmQR6F8ogpbycdssTvWGdQfB/wJ2dh6TKe+zykTqvOyWeTUjqUFQ8AyN
R1kT13h7T0gqyYLqNcTrOMgE6HG2hzxYmU0kA1MODp0RNbFC4EatmlHpuZeehBGSgMab1uB/IX+z
cbjyNJkGtwDKoq3F8nz8wH3abMR/n4oiNrCBkseTok2nDiUho1OqsfIEoGVI2rcMj+Vk3LT9uRkU
Q246fKQkeBgHgRRUTlXaa0RT5GH13LfRBcYQ5N1FNkcQRNAQgUJM3M6jp5ES8t+MJw6ZfA0OQfFQ
rAGlRiH1PrhjFr0bq0A0J/8TTqgrR1Sdq/yEmrr1cQBLp4PxNww1d/ENu9PHq19mx+wbPM35HSHZ
0SWpZfkk2SLm1thoyG8n9Fb5F0I6ee4VRFIN22d1xJZjzapKuGoFgNod6DYWHz1yZ1SyR+rthVvJ
f+h3aJ22gnjT5LjFDSCb6WPB3KC42vlyLuGtA/4ldVT0Zexav9eZM3lGOVKIli4nIiR3ixFMh5FS
6cqh8UqDvCaKO3W1/1pXD3/J5BznwJDwqPiMaOAiNCCQbZiZ/r+pHVPNzLxh/PjvV0vszcryBZKv
kQMfRnk8QBq8Jwq+GT8qAIk2FbDgsi04uY2pvCGNbe8XqP5bYS/eFKWymFDTMJozZyCEHUIVnw+U
ideIIpMyjq4316hB6y5uFj9dcE3/OUVL00x+0qePLFjQkYxn4a/oMzt/C5gh2Za/NOenSMuyRdPV
wEaCaYy9eD6POIP4W2s6RJt2guAFDamvrTD8obzVBifHwy54LorkqM1FJtOmCkV9dyXWBltretxS
5J7fwScTQOYFRz3SZg2xS3PJrukohA2zOTLAvM3OZBP8FDKr8EbpF5d4ZRF2l1zrhLoF9AOnWIu4
HQCtidLMO9tyszNijFis7V3JMbXy9ki1JTYvuliHeNg2ryBzFLEC7J0sYBQhkhLmc2G7ibELlo5J
/nL3Caw9Ra3u85K10qFAVa31IfPvXrWWdBP2csPAI7H9KqBfxcAB1Nxpuz2X2UzH+qfVXD+n5nZB
ejl4bih/zwMmG0Yvo6mha9+1K8wt8hMTIE66+6lA/Tyv2qxXGjhRkiqkExEi1Dp7EZE5yUhkn2+D
X6cY/VXAR+Dg6YVvT+gHK7XxjFA8vnfoJQGathfUiBmEud3jQeII0OKUU3UxKSCRO3yJvRhvOWY3
tTdKrN5MwhDqz6s8b3mrfN7pSkwpXJzyeHniWDWMiR2KjWzK9P9/vn3WNOZF7/vY/xeUn4H75htk
jjfnLU83KHfxEsa15aAEjNPrNmgjue4D+o09nN21NOT5vPGk+fgya/qq0SIAp73AiTrJuD+0de7S
VOOL0VRBHIKIBbNYp1zCk5A7eRt+VKBimUCEk9cQPjMSV/ofojII9afWC8xhRIixFno+KUTQG4FL
7+uCrUDmfHeKdp9YmDx+PSQHHkDyVf/lcUH6YJPcgyHKllX2iJbj9faJZG7mxCMlI1BLM78+rffM
fBu+bwhqxOY4nKTZJWjmAc+DNBYKxFKLmI98guBWj47wBVNHypkWoK1EFQxNrZJdE+gR0jR0dOLJ
JS5cD8tz7FWdynq0UKoSKk2D26ts4qBj+kECy3rOuXFi0CyJKS20FVNsuPMfFFxTRVIYbAIFrxDz
cIeXF5Q+X2NrAURUG1cZFoL2TMIDe6UCc8qC2XYjh64xgOv3GbvILjh5kuYw/ylVQEgTxOpcdenr
RyjgXIdPJqdG6W9YzLqRKRsLphThWwWrXnMiI0cil/p3m4JEbNw87K1dxT15hC8mF5NtQ2goFx1r
KDcrgr0nHzXpjhWONkvwUYa7b0Z2RfaX2t/jJpA03/ey9Bns1047+2sFzkk/AfAiJKIDSxrgw0M8
fAv5DbaI7rH+fEwevWGyZqFHbqCQVR4kTrfyUZi3J8Y/lOaHlkldVvayfsbuI0xYLEyimbM5MM4j
WHZea3D0+0OfvAi9xFDEoJrpYShktIfOOM8Tq0FQ2wFWBbXGxVAhUFB02wKtH/p3YWiMPycTf3q3
CQSMMms+38YKqVU6YnOWy2vlBEiIMrfWyNeZkb5l1xMQ8F20aQRRanA6hQjvOb3z7ZJXix6xLSu2
lyUjQIFdevi7Qc8VHcT8iMYudj5++ujhOn3h5t1XCPk9aCEOIcmf2hGNDDENtAN1FB++g4Qd6qZF
LtPmCKdTuUwgVWyL6JCko+A/OLMAd6fTFRmY/b7TY7rlhZdX46yB/8TCmMhWJjSdk1AK1kFdYf07
AIkwN0eEM/jcntKT+VuFsAoS95LHKj5VzRaj6NMSuO14YF49UMYlRN7Uog9P2A86MpXChOGOABMl
adB/ERcx54isp5rHtD5rjmKbDqz24HNrU8hYa97nBAldLs0pV8q2aJXksQJaWTIClzYPqLMxLzUD
b5hf2uAwHcPPRVUcqVN7dC9vSY25+tgMvOMZc9oGzGF3s+e0Zw7ueA1iYlKx5mfrtNc3xEz381eG
IsT2+RM4/87mDz7QNOOR4D239bnZWm3WviJgvtA/2q3tvhnnNJJsAoAxJLtWk8YSwiZqgFvJlvrn
Npl6hgUS8CIOWw/W/eKbCsXqUC1OGf6Cgh1uTXYaI0o7ykGDtVY3hrdvoKmc+tu9AoZQrAA0FtG0
vE6nrTsWaqlIzZcX/Spr9/A/YoavORYPBlYnnBGN8xW8uKNNHpkbLSeL/SHywGt/GkL8odW79Ui8
Ib2DXn4uagjso8rv1DetgBlB1tJmz6gLEgt9BCuMuqVq86CraIyZsBT3T7zeOdBSW58Er89JfUq5
m+GCxLRxZN4UPHQnqGODOuTyyoVvd1c+T+lXydmYdVZKJyov3yMscCx6mkevlISJUbBD8x22MsQ+
jnD/WeLxPPJhrJsMNR7kzChoWFZtYQU+3yCqiECynNQAHr/rixPlNC3Pp099XvQmXn8XwJmLA/Gp
zbPacscwiMboAn6+niw/GksYm7nLjdCArCakxMKoJ4OMs/wHMRL1Tv3sS43u2+vwdR55ZU3hz0bK
IqyFTO69ii1NxoCll4aXuxscYCs71ecbqw+GwfJHwARZxAo8RTz7OC0yRaEdSdYZgE0L9b3SjQiL
EqpRBF7TGV0nGPS5nw/TyMBJmxph4PGkkTENcjYB+FDg0aodYxiXpNz8lADc5QTeAEzzzfZAcoUg
bHwoAK1eeIeEJ49G00aenxVaLO3ovw78GMjgbawnsi+g11lCVUCUQxAKR0/VKjZsnrCslHgi9rQC
QaU9onXM9uLDr5OR24uY96FvSpWihxuXFnr+87ZJorS/v9p+97VeP4EKp2jDSNPiJUfmy7WfNqhD
rzUcT36c4WQVR6AT6MuFZr1Fg+3G/bfK6aNe3Jvg6jhVDgiwOJCd+qd5u29S5vQpuUVsDx8se9ky
jOTK9dMPuBipfDZ0anUzpErnc7+9kcCoCseMzljMR7bdVJ4GCna8rTyM85F5fkPdg3eCOuGKMGyR
B2H+xbMqELsWmgYBWsEM3jm7vVSJlJOOvvgOeqXyP7CpTn5gv3+3LrFFyD2hQMrmEq66KQPVVNTL
LJVlVloHo5ZB8e7239qUUG8dzIabPLuXQC1XHDzwx8RpQEJexASHUCdSruhGeoMxgBx7gWxynt2y
Rf1KfqTWcbm6YD2gLkLXxqtUyrQx5JFcDK2eMY/dUzwvHx2qHGL4KgoJ0gJSEY0hT6blbty6ZpDE
Q3wLRFEs+QvopPCyWOPKidQMlkj2sfY9GTO+jZR/HuWSl2wVMiKyZwd7a6wFa0tkO0NunXQpyEXB
MFknNAJVxQiMCc4Ecna7Yajh3kTi68U7K7ntMWCzec7Ct1jTHziNaHPVjvtnF9/HlEAHjtAb2QGk
4xgJEQ50dW7vBaEKVkp/PGk+PalgPhXHT+rRcy9vSsrF37xMDu2puahy1/PgRUE6UyP8EwNmYTXP
/Ye38wvanC6xD0RB+4BBJ09HBIcQLnH7lRbJEEExEUpzYL0YK00DwJLL2b4Qv4sIv+PLOyj17afI
jq5cA4WeF5zUn7GeHXTjAYY7BsiE6k36GELdc+/Tz7P/peurpfXji6mI+YzxrhkW9oIUxJ0HFAo0
e59k2C7zYjMbZbjv13zojZsKLyhbyO41pMc6UqEG7VnxGKZTlqWbAguYDq7qVdAemn4y81epOOff
2vXBvIDq7v69jA/7R76s7gb2yx+1fMu1qp1SBDG5nCMn+GTSiz5/E/Ok2KtiXMLgV6MHzCvDu6wa
Qu/hybMBRt99IaZ4xauUWCNQM7wvTD9YQ5s/sssS8sJpbqjOs8EzubWO6/GInbszkM7zA3iQE+P+
cWKYLCHr+KkO8FBaZkoBZ8V6XFLwCeFgBRPZeNmDZNhNpjyFkmYPJB0wkguz3iJTISgPIY0WaWq/
50rI5Y3gab2As+9LhT7pGR9Bz3CKfDmRJXBMzxMNqTpK3afQ3QLhcon/BAXbAYangNGaTwCIgUoI
FKNQwC/a4u7aiQz9RHCDpnjigzE9h8SABfKE2oj3+qf/+nDgNpF10b79Uw5XenwQXtRYZfzpu1D6
E/iPp1a/Aed+c0rBKFe9kHc5SiSJcFOiqIvz5biJTp5JaTqMF0rdnQig3SLFQRZSY8M+cfEbd+st
KyaswurF2GOCgNkattHRobqfH29Y6RONknRz+0mfAu0z9VmDx4YqCfVU5zeqJAVmLYJI8AybX9Bb
uOdo5fWeDSB6vWkqSVvGt6aGKcWtYW+kQD1fgpvQwvLb3kJlZLz1HYgkEJPcQpfPwpZfri6LikcW
pe/T6/GOxKaJ3dMQ6NoRiGT/BrfdRr9Wu53SusMaarr7U9OCdKYIGAD6ADDJV59WwcRAeITeZk2B
nT7XInZkXQ5GSjGfYJD0ktrMqnR3gcxKsUd8i+HxUu0DwX7cWtk68b3xns1trvgHFI8+z7rGmgRS
Pmh+as+NsTSyb/MWVqD4LRhFixvoiU7BBTXVWXpl3fiFQKjjbfKdhlNAmsuZrjINnwEEX4efMGXM
JiSg2CNLKLFYBYlCrLIgoSa98cvl//BzdrTz6PR45d60zm0Rz1kHG2UIfsWKpIdFLYJxPDA6kd5V
xv3ovYq3vjKvNNjzBxseuLaXSOBO9TyEYtYuCTIjMhatyiJK7wlFxd1u3HSM4UmczfzvXvv5Nd34
WpbR4TcXWwHvtfSw5EqHRO8GrskCDJa7PJ84OWsPbnmC1vxX5n6q+fTojqujg4o+qcb+nyTZvMN/
Rn2p0POuJxzOMnHOEMwIjS4f6tviJLO0+N5hNE3ExYL6LSnaQ8BCd1RE37GwtkE+4uDzy3CtP1U9
xHW2/P4m11m1gluoQ4rw/2sVC3iGKB0AJ0HgvcGvjLKC7pcOUkPI/hFHSz4S4fKHT9ES/f2Kd8LQ
kLsS1FHGduEcgEkKbH1PUb7suFOaSSVBWda/9yuuPAEhB9BanH9YoJCaYCXB74/RSs/JHuO+hODg
rxy4GwN+4FZtDwuPYMH8jatdubnQSS/ZmgfmkH565HaVqhNz0FzzIvRHQU3wgVQ77ssonYIzdwf7
dUjDzOrB2wGtaGZcVeuvAzqI2SO2tammu9CnWGsOJ14s3nEtlmEhExJzT392JxPRWQ70cZWu/R7Y
Nc62bkQvJ23jcWdciiGndA0CVAxAwqbXZGI2r+vVik7k7jGB7uOv7uYgBWFFd9j8clVo7nkN7w/X
gJgaNZhl3Z8Swp7f/HYMCAW7LEi19X4sMaO4a9DSpwSvrqRyIv84ls3Xop2Gokyicy2YFYVYC584
UGXdYvtKGd0JBxQTCKzf+xnWjXjV6vnysu6QTmqdeKOMdoj54eNsJ7umvzGeZ9N5EcS0XiLmeLno
gW1mLcqzZxGpv1U71dII9dY1J8oJ34kqS3CQ3ZDVo9uXvhfofo3Xn5T3/3S67LOzgkfg6bOcfKlv
68j2b3YN5XUHVPxqkUYW+KEmjPKD0EmR6BZ7laRWA8fZ5sCBL5x5Z60nCWhWa74rbC+ZRwy5a9Kl
tbI5Ps/xug0YfiSGcNmPcuW8PBc8euzGku4hYcOoGqyPyGjKx43586iQrhAMLleta85GMs4EO+Xi
xqT4P8PZgN/gGSFLKTn5F7E76oU7hTJBmJUuX58dJPEbbWx3xs4K2bwZbmJLH2MSKfPbDqNiNSCL
dysOI+siLDMzhO9Zh11CyfNQHK/+xNvm08dXN59QHB54ui0dNBtnEJ2t9lhwY5OlKQep0x7oPRgL
K+YJS5YvpOZnEqBZyxiX1ztZ7wZSUywq19A8Jnu0Rn3aYWSQy94dBU+P82zUqMk97iTvUkrrodLe
+79kEhE45JxjD3eZSuzVwSzSMhL4eh7yCI1Smgjfh8Ip0ugUtTrjaLqMe/4ssYCcw85Dh60uaBkb
uHgh/ryMKLiNxzSc7K2YZAhv2XwSkqjTlAx0+xxmh1QlqbKOQ3GbYnPLJNhRJ7nIBtUviB52vUa9
YL8i45lZbVdlDt6e3Rwy9pIsZZn8VJIyJtvGuAZ2Q/Zr9prCxxI7AgT7NjA5qwPf8LeI4D5ivMUo
j3tPQkePYq7tX6rsh85MNmzN2BNpY/4pQlDMlBCte4jojBD1/8h5g6dOXhaQX+tq9wqNoCcvJoUa
tbT+sWTx9oQXtHnGAm9sW9wg4ZgtoZ9FLbcCyJ3/9Jfg91yk5KkJQsqsQqZ0V+IFimWTNjhKj/nX
NiLj/inmO1gHbjL+j69Drea7QAKSTehJXykK0nPoTQuVwWCaAe7/Jbe1feMm8The7RP2bObCiUy+
thhTkYN2+CZpqfbIkCaH1bceTdLq2N/LKCLkcqoUmXbtunqzIdO8bwYDo922uKA8hHrCoaC2hTJT
BOOorN9mpu/0vUvh1/DjpsJbiEOK3HX/2V7XI06S5q8aSVWGw4jQo8TZnsIHAQSH6NJJmvUbQCuM
6I9k0xc5X9Rzmg6LIUzLD7nR4F1aIEylHrWcteVPvaQlFIxL6GWXXG1Xw4nKSrjhoiIlwtwweNP3
eYMw59ymiGmf39Mm9i3JnyolP41PfmiNva3TUie/yIT62p7OFAePurdNIjOyPrqH1On43wEXeGAz
ZbqMrjxDWWqL+tyyKNJFTpetpfOkqT5C5NwaotewGkOZf1bWNC4a2DVYXQCQpZWfVC1mKLRAnXHC
wWlfO7Emsw38Cvjs9eIg6bphH4suoijHz1e/PeOJfOnBWN35f2bJwdEzaEILfJsk5HNqCSWHHitG
OyR+63nTZ4GMhuFKsMQ3bdziGfO7qvXQib7jnaDDevsJUkKtcDCttp9j4TK7itYYjQ1ijQhSpkib
KZssOnLOHZgKBt1IYLNL0ymcVjdWUxrBlqE6Q8h6yz/hNpI71lZZnwPPKvpVdmAbwc51HpNPjmxE
7xnELVxdnCM86ASg8HXDy8lUoQHy9f8OWlY8FkXYMW0/5deRFBEC6dFC7rgz/kT45Z5QnVFMW3Lx
lHFLADIMNizEpbb9KpQe62KwKopmpuX+BS17GaKzOM9cbokP4eStrYlBFATNidJ8O0OL3N9HFauN
4cJYCEwPhMJ666OQKKMbXj8Hl6wi2sD+ve+OdE2K+vrpe2aWzvY54W/vzrrsx/yf08AlmCPrDodq
e2tqX6JgfzUfCRV2AGuRp3b8tiZvgwuCd0jpFRoxWND24bb9oKdQdBfDv2pss+aSKI+MeZM/4NDB
/gfYPeIeszLxfD4yQrFs/laqlReQQtYa0d7altjBScv9czZElVQQP6vSk0gFSkpfPMiQFwd6G7Ex
XtbLAwfoi03ZqVFPb05EoPXf4UruJHQtHLUk/SNMoxUnyCXulBkYswn2frNy6BmsCtw8QOzgtR5J
z8AqUKTD/TGYY/NZmuj1HZItqWQCM7/pVj/18TXi7RgE1jowrb/Z+A3vnM7vGBBhqG31ZyV4yjBt
F0TV1io6InmZiTqNX89UBRU1AflDoNxjI6AO7qPT/dV2QRuO1UKl+IaImGCbLTtk2LEI44wKcCsJ
miVgYVzeCyvpaW43fx8eAqdHUVeOwM6IzN0hN83WBe3RD7S/jdwst8fD0wVpGPOqMeZ9JpjdJqKd
r7RTumMSy4QsUdpY9A+8eh93nrd7UJXJKZwuHHXXsMxv3RbtXMPEcBv/9xgiry7a2TnN7fqOglAS
5690DtpSWgO2VuHBFwWeWo5yg+NjDJHithjeSUhJgcFS0eoFWbzV9GcBttP0gh1iJF4ff38MtSX4
i5NEIIFaSo1fNQysbpt83xS1AaI5uB82I11iFlwxswuohxWEGE9IOFm5L6rqv2+YOXpLOQ7RrTKs
v1uO35Nzly5WRcgFZBQuyJldhONEWpcMbdu8DVHgP49tqGGVLncAQ6OAhUvU1UUX6fQodeV9Cir3
9uitpWWeJWtAezoRXGaZW2stWTz3uPgWLCUVXa3ydMqs8yZVdoAwtCssTfriipTpOAUTH2PDxuJb
YCDoAy8F96HHvIYU+X1tguie9+cno4pEwlBbRg6F1vX1TUHe2qLh2VxA2WRsmE9CWuJXEPuzLYu8
RUn4O7DfZK2RhedGh+cU/E4adxLvkochSUFX8afQmacZbU0XscZ46TKHgIzko4ZUGRrtHVSDhecg
Td85ulyBGLhDG6EigtH2gDL+2IR3ufJTjODJWD+MwaNvpJklmN5L0nZBccD6KCG1jUboPDvXOzWI
X165RbIF1HXNHI9mgMXPkAyCps7ljv7ppC5gVy5A+PSqyJSPtIqNDxIvgtngCLHxTGUDHwkH1cPQ
ey5Xn16lTz/4fIxy5sdnKTzB1ruSjZX/Me5+fjiHMftML4hNDRcSzYrTaMwonxdlcPGPNbexxgsU
co35LqxkBMn5/LGwbSXf7UAH+2nTi5brSzfhCSpX/L0RFBFOFuqZR9wuoJaOIAA6YZKk2DoQulnS
W3nbzvgJFnaqazUCAcYcc9hUIiZeBFuvgSSbLPx+3VMesD5vZ0ITwutUdxbXPFmoEkFlq1hp20yH
ZW9BGNAjuzGbp8iqoU/yTap6ClLvh5CuasyK0mISwtPYrUxvcxySC4R4SK92QhwkOY4/3RAe9T68
W/Gkyzby91rJhaEvr15a+30zXXGRXYg5IPn7l043kLvaWuXywBXisZj1PiqjhXEfxt1UXRTHH/3F
JmPyB5CoZYwsP9UflqeTajMDU81/6YcL132HSq3iAuTNY+0V2NEd7nFfZ5ig5gbuePDsRNmIm7Zf
IzEaJyK/ayvEwZ+PpEod1Uh3ZoEsHJBDMQaz7BFjpVK7XtE82RvKqXypoQquTX7Oxe4R+68F72kN
65+6q82etWJw/hxi/i3VijoAPM+736cznjtFMWMZlxklD7ATbkgGakaBuM9MUctbFO26c+OrFR3P
aYxxrD2RSnb1IpjxA1hMHXm2w3BI+30RHBtZFtwSpDy2emul8vh8EzFsWZsOEUYuCzVk0I/ck+3y
lK/DAGy6aUYMWj1f+VWS229OjI3zPdp9U1LkZS79n2U9INZC3DNFHa/+aqXjDQBHZLG7LoSyshPg
sxJxC7sjLz72eM0/EnXT6qisJ5IOyZ1iRSD0Wv07FkpqcMsDHJ0SWF+Xo31VNMOOXYGcj/pL5Rxk
xfu+dqfWT3uBgfXgJ6A52DjvCcSango8Ztz9RZo1JpFOptRSm7Jdweph9jRuM2/5aFBdWZmy5GM5
s/kg7tJMIBbPbTptru/6ug8nNFUp5jzoEkQgr1q422dpcZUnCqInGKE0ciIwtCepxas6xOiSprm/
EHc42bHz/STmwfxVbOTB1CAZjbJAgSJPiPmx0WIBTGzChbUyQ+v3PDlENqKT+VjBLndTQPiqrF0b
psC7NUG6X62LJKG+fAJBG9lM5NLtsrsRsCYSgOHPwqNhBE0FKXEUO/cyxF10pJ6klEiZpMpusGNB
ccrfifY/5FVxfix9lox0I/wmQGdtrEUh9GdoziLiZtPTetHl4WmJPh94dxgk1IWwIK/V7yNZyzvZ
Rph6aJnY8ZqO1q3VCVWBI245F8JiWKptdtZVQwiFsAqhu7QDN/FohKfPgDsbsOaotNMXM/L0wB0X
vOfPQXwSxIbvvgAHVuVU6sylnl3X73Cs9ghbWROnMgKArniPd4zhc+H8wXqFfhEhcm55d6KmbFbL
JIy5tnRYDImH7Rw0SuSDPm9vpOCoYbD98IXjl8PVCZfBwgcMlw0h0U54Edv1Kz4/Z+djsSg3uPPm
wn0WEgmEn2O0xolgjYhJ8N3GRh40BXqXrpt0v1CHU+vAtliXut5IJr5hxKEecTaC+rNpn4I1Gdp6
93MxLxPYl00OkSXBJb57RUkZO0TEQOG+mCouv9tTPsbxIyaGDEie090NcNIzz2nOjrSN2Vek/LbN
xyptRuwT6qzgn7i4rWet+MZg6rA3uoFFsa4dyiP/pcA6sutOrrlMnaFpU9WX2QjJbE2sxl+Vb+SA
QbTy/cz0rZt+8itW19ZuSoITRlrMGOowY786/ArwrNjmBYBDd9plO55HeV3wgU2sB2uq9iO9Y87+
z0DOu0BkV1kIAWJVd/kJZXs7b2p5ijdamog0lsgeZgcE0xB9LMlDzu8GA7hDJdXbraxMltYmFc9F
2x1i1cHHHwyfvU+cjgakzMeLiUtV53xZ5pKdOmn+2QEztXjMep94tEmKXsyeyXV5tjYv9nonAKJF
eDR//XE1flDzTTpuZqnmXNaKlCg4zqWdGP6PJD6VwKZw1GvsbgwJk4jVwpkQeXhzQyBTv7Iv0LTc
gPdnwdiKFQXzOedXOtZOTxpIMIY3gLGTA3rDeH5SBWY8bIkP0SfDAbnsQ7YSZ/91Z5g5pfrGAA5q
dlVdh6xgYpFtDl1SUMWC/TIioWzShrXPeE5R91ewml56viC+uAQbuYkCH6sPQ5odDxHliHfNMktm
qbgThsqjr5iJv9YjpyiOtqeLJhbXrn0aFlosPTbAwHXUqi1d/WSdKwjhyq29MGfWwtay/tzQ9PzK
EOc8VpF6nU/cZcpqMFP/RW8UQLuxuHGuQvF006TwgjCsPKyOJBlgrc5S5srMeNuCc+XJ7MdUnnsM
JNt1u6etCtbBVgmXEzshWNCJOeFPiRdm3dFErb40Amf7rhXwdbaBiWC0Y+aQGIm3XyWuefcSNgHx
3fyd426vdx9JVY4mFpb3aM8t0IzOh8epeUzTGLy8lBnstgdnO/WJgmZl1kmkCXHZCldms/ruMe7A
pcaaeFniqplJO1wcZj3DwHKUWB4PJioBDkRKzBFBjnq/t3uLPWw2r7HhVa1W81zm7pnMEv8IQS/l
gw2Zp8wiNokNV1ZxQNv6LxH/ndYIDZzB2wF61w336xnH+odvOyrxd75/QRcx40Jk2E65fUQxF4ye
qBmn8ajt+/6+FSg4KChVEg3Xx3ZG6lzMhGqgzoxInOCyxF+yXOvR8eHwOFSODya1/9XqV69gLDq1
YtzA0gOYYPfpi5hsknD61+0Zp3R8dFggJr4qY/Qdhue7XOUbAXNbtdVxELHBSrY0U9w0XPUSfCHJ
WkH25WcMnPTYDhM/+NZQg1/l5JSCNrum0fhBQqhiqL+0+WHBxFbYU70hrrn4WzRwbyr+oWEr2qub
FI7u+H/DtUiWUj5d0HnqKgLVsIJOmvuJebNvGAmtrlTjI298L3dJSbUjQRm1tslqGOwXQVYRkIEL
alrm61h0iFqwWR1ijQI4wXYukcfmiIjXnh2RnJY/5Tu5pR+AJ8xn1ULOlyLoM+C6YQn1vAT9qErj
EiFP45AgCrVuahs7y3biF8CrgPNi9z7shqgS0QbYW4u8uzFsuM9U5KyN1lQx8nnuX35gWO1pjc12
2c8l0coU9CODji+rvX4RS3FrWA9zKlo0uyP7UEVxJnnTUKnAp/qLlXITJTax6bJHb5nx0IOfqsVK
RJIuLs2fpbn6qDf+KLEt0NuAHD1WNXPHDbPGczjoLdj8jF++Cdg0KR5rM6lsx2dRy4B17P5ObuY3
Aq4eQ30jtToMHKrI/w6+Nip2tK05ET6ZTUdMEs6vcZZYb61wOLRs5w9lsQCNYj0OYgZCgBeL9p11
du+lwbXcHPb3Lsa3is0RftmbPhJpVOEhrLgFuZB2gVeHqtyOmwVY53wWmi7B8wijUXHql+Ri1/W5
XP7znnJBk9Jy9UqjSE+cxVQfC1SoW9uIu/a/dAMpupMP/4lAjUWN6AIQ6KyyxKWlFOb+zI1iDaW9
Meg1RpN/shpMjGCkOMxIGh36PrDRG+f+UZN+yw//iFKf9OK45oY8/5RaN5Ho4XHHPjLxS5E/k0Mj
Mo4cmDqclJaI1FYMLKjhRT4Xp2i4AWlOvP59xaa/7QcC+1fxU22DxX41EnwumZQwhIiUpMCUdru1
6qSozySJjS5rvRjhoM0bwyFY8v6BwoaMUzsdNF3nreNE5jP4Bp9UzwoMjM9nOhskaFXt6vI6we8n
ss8f139mfW78GMS/gXbm8A0EiXmMrR2yNOkppwZ0sBUVwXxLkAzU6N/Fwv9/1yizZo4U5KgsW2MP
XgisuSUJC1bHMU0uuYSNurWWZfTjOsqqvZ+yJxAxgGQySlc25GPvJa6LjZgZjbzt91bWEu26YRqt
JlmGI34in1K4luCbGqAKmStf2ycDlB1i+SHiH1NnE6usSx4XsJcHU2XoLvoLpgTOSDt9Eh7v5OPC
e7ecxYtWNnjKoxLyTU2Z7DntxGys0ucWpFJOavTryzeeFqUZxPIWMnq0vKd9aGd+kdeKC6Z0h27m
NM2hQQ1lYxjPZlaGNWXMtwbLPNfQm095ns1UaSYH1PrliviAB7rVNK1YPOOJ9xsQ4cL5C4UDU2C9
GKwh6FfH/uzr8KvQAEc3xCFf/fvbq70Kko4Q/YUXZctv2o/mU4sXb0COGECCnPkP6e2+yqqrjptr
SjOPEiTkTl4bSkWJjBeHZMUoEf1SefELpvJtoqdNx39IhFH4g0stOWcIXV3RHuKX3ladpsOU3fiU
+kJwH/4xaQoFfG7OucSMFmod4HBtUQrer2Ai8xtAfR0sN48IGVQjrZTnMC/lTpvOm2kk1d04a/A+
wa/9PTkmOYyhGyDdoCe2ypkZdfjXsea111C4s90XUvvIcR/lp+PjOEyINwdSj9kT5TxQZM0xrhRy
dkI7S8LEGhnkblYV92bGwaT3i0Vs4PQubyA7Xl8D08z/ZEVcTYZmbXCwxAnkto3pLMs1OWgY7Oli
cvKnGKL0Mrp4kwJvD0ubFWI9RMAIEFWvXT1kOsAOEykXSxrehvyAqk+nfGFUDSYHzAZ5BTSWkWzD
no+4MP7Bif6jen3/xPCbeu5SaZpmtQOG9kL1/BDiSK/pVUrtRZm78dx2HryiMNC08yOl2g+eg3nz
go5RNPYjwduVGTa2/y39JYTRjT50UCm0S1BIKJKr9EAZ4KrCfw6mQjJVblNtcpDRHvOqeMQJV2qA
cmvJ+TBGSwYwIG9v6J92diu7wukrWVS449Ei7HdodY/EWlq7x+W2ob/FJAoM7LD6Hw7u9tID71Jc
jMT8vJYpKsiokhRuZfEm7lLZDmNQwSsEg7/ojj8hMRkRm4UWlyjtyfz+huaBSMTWQvXkxEZg6JDD
x4IUTOnELhkXD+YvYYDVKxWCc7DxAxhHqBiSLmQt7TwtN5F6I6LECBWa+RPqpk+1qqvPEBcCKcW8
/mDzwBTLmEtqRIxr9K4gjtm3vmhx/KEmbH8U/s+d4oybnv9I5jsLqc2Lt3OSKBrjLcIk+IUNp7a3
aeId7Sn7Ex/sYN5D6ydfqLXBO6UttKQJSPz6CmeBVHWrMgTGRWn41l5bHuNGGy4emppTGpi7Wzj1
TUtViqgR0nbOliQ0eXewC2WtUe+dq1x7Jfn/Zg9su6ypxXi12KlqVFRzdeGbc+lJgYFMM3SUflSU
6xxElfeK1aOHseYbBSEhNmAGtOPlKpn64vcUU6cQzIjJRbpH5O4vgQJpWLjfo61nsK8lCoOwedqB
EOUuRxnznwe4TW8hHo16O+wQYT0FYxNJDMv8kWArfTSGZPqT3jGUtw8RTcpixhjKpdsWsgwO4ThX
fQEiUd0Pr6qI4Hn8o0BCwsxOmxMwaBXesSAnTx77fBRTqNN+bru8dn7NO1ajJysqzBSP4wB4Kob0
RPIVXEMMqxH7q33mC9XQ+YfvD8yOsuCJc/oE7EgTOdDUfU235tYOYW0Wrg9rnbRzYhIEB+XGnHZQ
IOBdOvhookHxcOtQt/4c1sfDMQxFtbieDwPd79HlVObtB9vnDk6Guhr7L2v1IP3diHVVWeZjOpvD
G56TZD98mQ4FNBIBkT1AFa2e4p/SLNed/IjqzPgheuFFd5/r2Y2l3V5L7pXbwjyEzmRHa+b3p2u3
CfhcivXPD9nHYUfo2lrUKu/lUR9CgSnVv+j90hIuj3I6TkHrCEk3lfZZ/gmdma5xGzHqWcjvDkuo
kVsgnvDL7AxjCyOjqU/oSZevEKn/Xnogy+jIDsUUfhZ33jamkTvMPCcYxmyrwy+4hLE/hQ3//zkc
76uKYd97dlAfUWk4hUF4/fIFHknDyXO8dNNOF2lBjnU29uKZCguC66S74RethkgVMU9c7wGnMJuw
YLKvpd6tWC8QKDbNiRhLP8tt781YB//XrjasqLr6jlSwmR729Aq92oTkFYFFFp7aOPt7Vtka5S6q
py7lFzLZDUSU/AoYjRDII/TPQmbgKEHjSOkFYLRmFrUvnvYLfnghWM5HqaNegEFsp3cAS3kVbcVM
vNDZy692ZTOmVoQsMBbmLUgZ6/AV6Z6+5BKNBbnOf0Z1+1U8pGm9z5Xx2B9ardGQ2hUjC2sdokeV
KnnQQnPBX/S9HJDPXOyobw1826KXeB/D4CITMImODRsfK4cBKQMzInkkGpfPz5U1Kt/RTT84A/zt
1XeAMOOXxyH7PH8shbRLR/7OBAKdHtD7q1UiPdDP6FvdMq9i8XuZuQXr8ll5nzXqCCYCKQP6JomB
h+w7MfQgKRu0h0UxqyGVsYm+cMWforYSvr5gc6GrdRSIq6Sb5KorM+SkRHcRK/N6R0JFp99R798y
pnE1OWSKMNdE2SKlVX2aqQ77BeWxnFDlZ/C83u1mRcnJ3xN6jHUfQkJ6KowfixhBBMXPmqsmyp5h
CNv0SVb7tQptf6GkJl6ouzvfmbED+ZYHlzmm+2Uk+VqQsv+mvHa0io4o4M7aeKGibegveBJpRt8+
huLjLBp5qpcXeGQvTghaBTXJmQGHT0FJZHoJyqXCJuttqEl+z0uBWDVcYsB+iXcUfn595vNGYMZ2
ZfE6oA2Pwi5KJkil6qaFsnyUcWIMj4D0EKVndJvBbWpKPRVSKasukAWteM28PIG6uyksECzfUNAl
Upar2F8K6suvd6EWDOl47r9dLXxaLQgav0g/zjw9x8VvcFBixZsOjXGl79s6+FMnrH98Jgv8R9Cm
bcHNEkV84DrcxouaXHccYniWHoCfw5chgLStiYII65epzgtl6mNGUPeuIhwjBqbtjYe/VcQwqrAA
8suEb23WrpsBcNnVcI2gV1aLp5UYnW9349eFbm6YB9CtGeZL+h/Zf9CtNAg8Y8/o9/m4NUi7AO05
sfm/YzKxr/+TiS3Ubc9UFLFu8FTfAuqaatsOrUf4/ohIBqLsBDTK3d7R2tixcnsgoC/bdXf+Hzq5
lhcyOhXq+Zt7f/p/0hYPpFYkt9OFgmfuTSB+upGDqTpAwzP+iTvsjrm7M28HmeDoXUq2nlXepMbI
7GWUKKrN05i50hpuinzl8TO6nEb2GWOmcjussGSgCfDEpeD9VDp70xsF2jK8yyMyuT/Ah3xS2xI9
HM7wkBEYrlQeOCl/zervCVJtGQ3Mll0txP55Mk0skpI0GCF5LB9aEsFGk1INKrQXEGAkguxKInyF
uPt3PBZA+mvYOMMkpxUaYqweb5vqrwRcjx2ZH9z1obzjcDbc7A8vFVBqa+bQgO/BrWhSZJvWpYVo
Ozzflju+IRmOhAg7S76mfBuRZ2tVpNX0tzIxwwEmUVhl5FKvVhgHf5gAor/PyT6A/qB/huOIawfI
9H3HUa9LsAYIiaY66rh3qylyM2lK6JcFwHJcg2xNtkX90hB+69EdV5yp652U9Pg4A+ETRpoikm8t
Pe7h4Y3PV0G8uzkoxmTi87Z68LS3oq4qsP0C0KWuD2391wLvCdBE/ev8E1ZRSBX9MGmboT0x79WB
qfszLnB+AGu+RINFRKg5eAXx7IXc9IQDbLbNDt9GLtuEzQtub0hXL+o0nPkckW5lKDL9pjyUEyAC
N+jNjaWGyqyIU86Bb7nWfM2oTou1hSBnzU/jGe19J/bjMZXPx/JA54Bu8X3szmz5qsCGkNSQZKZZ
ldEcXL3/VUmWC8UX6zg5kXauXrRFlo/+l6y9Arja/U+smXFhsircLobgkar6C4r3rd6+8jeJrru/
+VoiEQDZo0c89vK4AOHMePdD4lS7orm0aXR2j+KntLTpxcm7y9zBc+uEAWl8NrPrLzCk26exNMWa
q8V00zOX122KR4iXQH/R/WlHveehWm5kIY9I9Gu46VrwOvuX36z/IiT/dqOg7VNN806oDUtzQ6tD
Fg944dIPHuTLSdUXLFV6PU3/ecaXvqHw0NYsb6dxX4E8QEcmleBZ7c11LAqQuHdvqe7cW9nEpWsB
D3pO3uBgvjVESUPSiaeQlmZMTk1BKNrOjfn+NyMBy4q5b49T+d7wjKY0rpDSaPfI4USY2X4xVc5E
aBs20GMm3AMK4dcn1U6sk5oNP7lyYtlAhnzfR0s+q0JZkfttwgfdw5vJi1jMBcS5cI1isGlHUBYo
jL/Hi/tQWUsHQWtVlyEAWPJBwwAqml2YlRNTRA2aiRS3FVZJK0YOYRqTIGJkiNnLoYTlQgFXTJ4i
NnFhbplNYryWug+2f4kuaKy+w3e38HYUYHnlN5SpeAGiVV8KsZ8H3uVyf4thFRracuPfyRitDKC0
OrWruPvvWT/tmBshAtgRdRQpjekistLmKjpfYFpW1I78nO2svAFpr87KgYEfayAjrMr+mKaQKvIc
DaL6goqkkTJaPkEuxGok42gaQgnpErF9+qxyjecmXqZMnjl8OV+VMuF87eUqYCTfh9Xj0i3SEEZ9
Yq5DCRuNAIcsWnhBaf+S8B3rLm6+Ui7Ahujhz669E028YKk0LgNkGtxax9S5qzrPbuniH3lHA5Rw
uJ4Uw8rzct5NF4txH9mxTExntoEI1ZcG7NqtG/ZIsJpDbh4/wHyCnFVXwpzrxEPOVrFPqZHsGBil
x2F/yfrxnuwBVWRUkcSQpUP2b939Ute8Hp9ueZ1XyV5vmADNn4SZsqT0atrjSe2EZQjCxb+OXY1/
ODsHadcVpqUW5NragmJST5C/PDIdcdnXxJiM3nlc/1jGI2fz30a1gwC5KLSLn/VFwZ5fGgCNWobQ
3WVTCYbND51yS1joCxMFZ4xfEqI/2t5gkqmgwkpUZgp1vjHHQnZpVnHt8MfSGkNXyCX54ULwv+y8
IDJrBQqJ5LnyX+VrvkyNxUO28l1gHR5VBZ/2CLUDpV6yHC7PEPYnUjwUFiZdWetbL0+xJ6J/1pac
zEp2iCy3GunclQDD27mJMDWJI37+k2vauEIJ6eUYGQJ+1sqsAdoh9Gnwu8WLbzD0AuPTiNrS9NHW
5hNc3Yn19J3YYslywtYNYOBq3yPzt8rFWTWRr+GgJjq8oS9UO4g7hdmnR0b+RqTZ+mG6/ZrNLY6F
4UQtKgCkOwWvC3toe3n5i/AwhQXUIIS5XLZMEqya3M07n2tLHd2Bn1n9zWo260IJme1ikcn5Hv2V
hgnrH3ChVb89JjRFKWMWuMv/GOviC2UQ5jXTlMwMrS0fsig6PCudHihka0X+qLmRSPFJV3U9hD36
IU6reBqfPmiLfytEntCh0gJ84lzoJtZQB1MrJdTvHfQC+jLjflHDtU3zbMMn8AdlNrNu5AbtbXlv
yX9M5hFmd/nbUqubNHz4Vqi3s1ycP5mWMlnrCxJSyRvKo5XkKaQGXCFs/bHY/+xCjubLkpDeWfgI
gEs9ZD6PuSrOcpAr1eNYHZu/raGBHa2Vuh561GBKTps3/Dmv5+12Xa5UGujGAGtY/1MP/wlLHD6y
n+PLWDHFX/dQECAJE3nbL7eHjhW0FzJrnpT6Np2k80HcGiC5MBnOzOGgo309m09zlHB+ul+C282v
2pepkDtxp71O/8nxrULqWqPpXagaBlJDE52hbcRN8eL14TuvAJDSpEgZZ/XFA/1wE9s2tdNoOu37
W0SLjJO4UvccucvfIQCkp7x379excCcw1JuwPpzNcQCyW7SzBwAS02FpkbXonPAgbk65GvZpid7R
fomNXOKbrRvyANG8/DN2NwWlenOCBxEN7RUvPPcQaIl54c7prcvjOVTzEl39i6XeIsOMqurWC+MP
k7R7FeIz3I6f4AziOoMP/MjRJlkJWBm62MuzQfu7B/rzrvCl8bTYvyGKDx0anrHAa2eswqQsSW9E
FBRrdUEnE0O9iQdwaOmt2xX+uJEvI0lD2y76WsDXfLY4U66hUhXST03S7Nq3MsYQv441udHdrSSg
xJAD30Q1fzP6eLBu30K7hP5dDdnFFQ+vpSlZc0n2oengpnUHbtYo0HRj/kU0yc6KxPwqqU6KeiSQ
9h2QQV4Xct0EFvdy+a9byZDOcH2Q752Hnkxl6Co1MOT6rBw4FFWCyl0AN5HdG/v4FCWvnMAoJOyb
P5RJDpOxFWz2LaAtcMFag7xrbCKoI2dPqdfbrvxnDoOdphjhz2kdjgsdrU4+FFFDDbWfCkfN7g9B
6GRpsYVXOZzZrlKPYrgWLmaK3cSvRh1rRdmfXaKYKF6lroxD0Nik67ic9iTOBLY1bIPbw+LQ60IM
Ly/quyohuNLEWlOAVpjnidO/YcwI8gfM3zdYhGFVBoP2xQj3wslqp8T1xKUGCGf7UdgQ1/7HEY/h
uzb6NN1sYz3dwJowTYERsIA2jwLwstGaofvSqCx4t2clS3ZXJP/XXr6C8Rd64CfBvkLsElCPWMo4
AHy4IQXKDxYRarObxkupSGRPi+uRE+a20LzgF/y4RUx60jLgkcy7klPDSx2oTPwin4k/iCFdRlwV
oD8wkZR5gi/+m8mk/VtokM9jnBWm06G7fVb1KSsRwDjzMF7i+rUYeqon+rLrqPhjmYAhtjBcpQo/
cPXYzKWZvZmLUJpIEkcVCyMfnwaz3MlQGj8VpcBSduTOKeadJUELwO9rdtT4z0CquK3Zc/vipJ1+
zzTNxxlmX6up8qJarAgBH/76CpBRwl5q2n9O+yV+YLOnGBUs+VF20g2ooIV7j4rrFrwFfVqvU8Wq
sOh4ECS0iXvpFbj3JUxzCSYDcoa/65C9A4WskoLiEOD+Jj391XhnBNl6/RltOubuMu/EBMWkKaK0
1j+CqHZPX0TVeYGis7axmb75KOLM4T1fdA9i6qLyNM27XwW3aL4TPAkppV/SVDawJeRqifvlgCGY
gPWWtaQezTXddHBpS0BLW49Ge5+BJevywzohdKIss+87M9Ff1vJpCW5JyQM6TtdNXjPnYXFkBWo4
OAAmInD28VeRTAgclNJR3ytWNfDyWC0mn9oz4lLuS9enbkhx0G8sG0Djg0X+zB8JFDLUJEM8SxmL
qQN+sPx/lNgTTrjhZYI28aWgxj1GmX0bUtL1x7VeldRZzlToVVnyvL2oKpigy1Oa7czy8ionlX2w
OX2PqMIyd7FtugqdbGdSAz2ADT1szW/XlIjLmeuK8Py/uBQqfPjGYbLB7CHNKxPq5Brj6+zFqMG9
irSdn5f92vNKPN4EBVdLcvGAyf80RViv8pI8Wss6PsdCukzbfKyaBQ3bC90r9z1yBrunuewkJf1M
DvgulUGimS0RsKNrZmRRIpVgbpgL9Ctdma5nPSF1bzirNnkb8ZO/mfbqN3dpDKnsFP7kiPhPK6oP
n/H1ZRDuWP2FaFoCX8tverlPIGnuPv7TudOrs/vjxjw2N3bl9vCE2VELkBRpZsRfkh8M9ZriV4SC
zgoSOVKFGYyyCHb11XttTrLF7qG/zBN1DPeeK0CxFOAQFE1xphGogBavQB+FqzXYICQnneqyyqEz
gm6ugwTb86tIfPvQbvQUF5ePB1e2dLZ9IYxkt/NAMU+sjBwr42FvewpeRwh6KogEK+MlYKiXA6bl
laXvYoypO2lWSat9NZQXZABuEMVj6hSwSp7SIvbhbVqrjfvqUZ+0TbtGuJm+x5bax7Gw62RWfVXn
4cUaARDn8FNSZ7cDP0Dyz+Lmy9+DkWpL1TkEBr07Mkf8esoFNxvL51J/DYpjvXO4GsuRLvUkfDmp
IoxT3KHlvaJspO/2lb4JD21EZOCyGkNOU4rN3+lL8SY3EuadodfS5EnhTwyJ622myiYhvWHOeUXy
rHvRYNEfneuauOzsHXr/73XAxXRcFFM9LmiXhDF7JQN2mVPYG5D9kt1tPYpLlIHBVVwLOd/DyrUx
RF9ep28kIkPc4AblXRjWR8VdI3QPNyuANHDIktY7jYGYYos3Tfc97RlUthedT3vaHku8wxEpS8nO
1UI5qon79J9ll5WcOl52j220wodHddTESIRO/wRbnHK7QjIpZKq/TjJf4Prmf2IPRy+3Kn8B3vFV
eAvHE/f50Niw7AeDYHqcKvWZQ7iVtV13+e+oqvYY+Foog2tYjkwwWwbCD3AkUCoMBe9/Q8kO6lGd
B29ynLkNTk+J/hIgpgbhCHprz/xBljG6ds0N4jW1j0gxUd5E3xjQtD4bX/3b6bzN7P1o7xHNJOee
vsrzAqLFB76DhQTWlAmfHTgVNA0pBvrsHh9opRxvGkqU3Ra0U0zFbpQk2loTOsF+msC7G4BKEt0c
qWv6wUSIIhrz7AAJMhpsAUQSBxmiJV0f+LwlTG3UyEwocrAiu1+purA5FKKEM/KUsNuKVwjvNAMP
Gph+WfHWxALmSwABJ9hkkzOJYI8Bla2vu4oZjEeigOjrVWVVp9hbkuuCk+DAlfcG35ZVsZ33KrmL
nEZDpXgipcE4LyatKGfejf+kKewlBPDqtJMG5CTaX/1lP+1Zj8pHA4yT/qv1oOdjWcLHkAR9lIpT
mf/2BD1maQgHFE0h8yZhJOvIknygj/JSuzlgiZOD/AanbXiOWcemhLjiYfZ6VkcFJ/umB3q0XYWn
wL5g5l6sujLxz/8KF90VlohvzcUSrZMp0phLlrgLKke8FJKNyyGFHl+92RSfcKJq4vpmGKwEHMux
bhhjU8+li6LaNxLlMs8Mx2SGTb2Zl6dkPMhdrcqd0HZ5gohXXqURxQg0zG00/5HMKgTvwV4Q0Bht
5NFJuj2uC3lAtf+zmgufHop3vQGbbItuJJe86OyYx1JUIIyOU67c13G3EHUAk4HXMJLq7diV2ol8
FA3gWxE4hXBUnUilWaNkO70n8MDjdtrvw6NDEybAw8S9GJ8gQol9px85T2huOvPzYIeeZeufke0x
uEEfi2NVAlX0ygq6VuHB1h68TtHT4vMF3IE4nXDbdfOO0RH1YcUMeMO53FtYA4Q3gwieu3cr6las
bQLka9wQm8hZ0U3pUBbePqxCFgCsDbuX8NXUL5pDTK0DEgxagK3xCU9cfeWD8DxGStuEqERILdJK
dmakkKSsV94kKilfvD4VbjJizMxh/Adn2JAHevZrzwYZZ+Ckbss9L6rPZCqgOvTEpXFs6fxbv7Y/
PXc2L8Wt0iF1P/qdqq8QQUmJQ4DXcVMJwRVmE5HgkvvdDrF4OhKoTRZvV6SEv2jGfpjSDe5XBJDu
a1zZAuH6gAha2b4CghH0LTspvebdPv7BV8/K3QuXW7VUB9Vlodx7UvgnwaDI0PTnR7lcg/WJdkjj
RjregSfPULZ4KtpviM4s6lI3H5sqc6COoiec21P9spQToI6pnlQ0f7dcyu7Bfo5JjvGbUiDeYz19
C56KONFcTH7se6tSEB/F1vsUSl0laZGpm/HaGZ3Dk/IO0bqNJuwZJjzjAf9Sl9H3sa8poP5UPvdG
KVi84evDthRAefYzC8EbS+HVULSmAvbK1Lg9bl3X3hlwf0ppfcXjt19uI1Q+4oed202EN//Ineji
gH7NoJKXyxfoCuUqd3AIJlUYWeabJUxzmMs6QQadY0XO+ph4Mxr1lrHege8PEpTmR7AYvVlpFC0z
DKzOKJz7+6D4ahwaNnGsayw5txvoJzfSUiYqukoVrRmwB+/9t6m9Xe7Mzq5B9pZEYQUObra7/qIR
+0URBER3+LaDP/V4n7snxxDIgHeSJ4TQa+AIBw57onI9lMe10f7He66PeDXTConW5A2XH5WPtR+P
psrJusfvYOKCQ/hsXVp/zhMGdhxUz3Y+N/2dpeaw+U1m4v/pzDpO9T/17LeoaaDtn/WMHOIqwdCs
Ac3/kgfWORytbxD+viE3bmpP41iet+hAFPhxZbLpDcFBCcOR7dNQuo51UY58TdmH0FHBcBdGbGhz
2DZJOPmv+tAuy95bqmVIa5x3yxswEO7bDifHC26BJMA4NUpvb1vpxvFvvMEii2iNVBauSIY2VsmP
lhSgJINhCulIxSkGopGqPnUA2iMoCf+bLfakRSYJSj+5P/AKgPUarhZPRw87ycajVupvFZStVupe
1S1G1qIZQOyEnZWoe7On5MtxjE+tk+Pl+P+A2fBJJpIXipRMJruogVouV78qblMr+efMppe68DVZ
NCrVyZBbIF5db8tVl4tSw24DuFPTlqCFuaaCJ35TXeRa7dYP8vmzkuxmyaRv9cukSAafQM7VXJoH
IgAAVDCuKqzs+2VZuIsItvK973E8eWMylkWAFgRHvBc/P0IOrmyAtMQrUkmUliXibslKUFpbCIrb
ay36Z2qO8tBaQu7oapsDw8qGvU3+b9lBFYKK6FXTEJ9Ubwh12hplUVhudoMlPviiw7wnmL1uZg07
EVQewrGrVQnf1PSra5kuZHcT1ezmiy+CZJaUZgbHk9RSbCsGiyyPJIcm+eRp7ZhGElHwDzs0WvJ2
lqJJ8It8bdDvKwzarm2eK1UIs1AiUghhaIKVRahcSd9+AH9dv99iogfwiCcB/2DGtyX8pqI6cHEa
XZYyV8h8THe3ffl9retN+GTAdd+r8zeSYXKcblWztSqRYa77Nd+G97o9JxtclFVwX3W456di6WlD
9Ue3j1lj8pP8meF9kyG+fLvbHAwK4v87ojNCmhZ25auHEPtDOqNBhEsbgxlIhJWCsfO898Pnyavd
yYUaLCf02dmmhZJKLKRfDOOtDXEYCg9OejjzKCqJso37KmBm8j95j7CPHG5iOQnbFROolFoOpm9G
GaMGtlerlDcgdM0yYazfcsidsODiOAInfwhJTKmWO9UyLsJKtCDDary6WtanuaSpbdEiS4z8Lxyn
kOOAH0kJ/CQ8V2V4RVMS/hUP2gdr17Ptzf6BdB8B6mqEJq2drCE1kuzPik5CRWI4ewhCQofDcPE6
1s9wp44wyhlh0/4ne8xVxdqHYobRsVgi60pPQ6s8BCIkJtfYd+fTQuyB2BHi4G6VmtGfuH+YuCi9
3yRqQZr63dh/E+35+pnw0wk1F4iqciwPFCW0E0+5xlay7bazRrkB108JfuBubtC0avQhBqxfvrXp
4yI9dFC7pVOi0GSiEhgYb2HBu9kSTKiCs9UvrxwYYIsbzKvXoyQfLnDLDCOXmIToGw+BVxjJUknA
8uKC1A1Rh/qL8jtDKOpI99fyr8xVVtVj5sI1ROuDm7QQUazxCeipNGSf7e+7fbOktHIyP36b1D8m
KgEhLIxx0I50H9iGQh30HYrMted+PDPbkYu2ka2AgFdr1j5dXAcJGjBaW3CCe7HrClG8Qf8lSI9D
bSF9ASpihXJ7ZO41/ap5T87P7DDPydEWZmvlsIUgsbbVHS4EcMw97bOY+aXfwkh37C2x895B5Chx
sDYohYFiajewheM71B9uPsYgdGIolaME2hm/UjtTcdDFKDLIovjdlR8XEqtd6fO/rBRtmAO5tZwQ
yGGuebdGjQ+6ZdKeMsX/4nHS4KrnEzLttixsqgS/kiJWgtN/H278Kagr6BI2FoQWpNLPO4lvnZTA
eTzMSfeHC1A62xhgdXKVnY5/f6dxGrRElvecmkJeRr7o2KIYbH+Gg+Jys8812WK/z7aXmw7+FhGs
BKtY2QYQqwCzs5qJ3s3B4Y/XrYhD6AF8pwlLjAMGxhzxl2lSatsGTnMoGA0ApG0h+g3lgZxipRk3
Cq+Hx92d/RTJWeE8do5gYQzDkbiPDTZ3B9i123Vg42drHa784W0366onFrVLufIQjKgjQyVcNL7F
9P7eQIykq1i5LVkqFPKp7Ma7f8MiJIb4kx9oy7gTkD0jJe2DIUp0hTbIUcRe8d/IbC4XPrv7FEo0
MTXUT5+k8edFGn1dGP6IxjFa1M4FNsTunaGInoST0PSGn8yJ2D7dKJppWwUpNjlWjYWjkXtRJKOA
6kz8RkkXosB5w0l5CyVfbZHpZapehcQX0n57v+yXzvs35FbXVC/T4JaYDudvHHhjfwrSBCg9UXLk
hpTDKnZ07vcKf5elNDqWbxIlCK/jXMZqp+ado29BRB4+OPSBNFVbjYgW8UwueGLGKLf7IWa00acy
ihZteori41EGeG2bzJSWe50J/tKcS0VC9Wc8KW4RIASUxLXaRHcaFcStbhcTRAqmrnBOZ37WocRN
TU56uWSVOR4PedEJdtx24BgzLf7ASqe19EAEDrJeG+gWmKEUDfS0vL38G4mZBR8OFm2cAMIHAdPo
QMCa+cYnsZ8/VVFlMsbxp1YT9OWZ5xSFFpqJzslRo2YsfWJJrnn3WkQK4d7lL9QVaP4jDcSM8wnV
K959sWb1otJioQATlhjJe232z0Y1+7Vhvb6jJ9ikVSd3onlb80TDMOu1AkbTots6G6mo1E6UWDjw
/kNpeeGQjcmWMir5jLB9EfrOuWXsTRdPmGtCgp7g1BTiWB4J3hB9lqeXEXlfQ3mgX9S0YhztsZ1Y
I8FXcG9Qr0qWPw7nlzgCTS1Vy1jbb/g9cCZDCR5aN2IirG1hz74+PoUp0WWG4ebz+9K10TYaRSVj
v5gmuFsQ5/nJF2yh1BKkx430CrL9fFGlad1N9O8tH+Ubkk76acvgvz174PZX0xx4eVG18Sg4X6Ux
bV/dYXO431serQzJMle9K97ZareKMAln8x8tatWCd9SA+sJRDf2DyyTcpUwCk/+Bci+tAEpx6XZL
MxKMN8X9cULIL0L2IafDBMF7RX1cdhplRL6sv6e3i3Qv81rEFStUX/hLsjYpNTo17QYSM7aaNl26
AhtbIjy+9jIT+TuI8hU3+Z5nXITRQ85R0ceI2iKjJ1Q4PAq/KSJDDewIlV8bwJctLAUaf3ka7ouD
oKajFj9BpeTaj/cYxKlwqcx7ljrm6U/Ujzs9D/l9c+4BlL7NCg6cxmCF7A3IdWCkNlCm9VSSD30r
fPz1ZTiqoiscJqO7ylu6Ts+yTesErgXsrGgs1/7PPlXl7sOrf3djTGmg8ZF3aCfOiUi0M2kGwhsH
uYMqTHxO+goezwo2q7WTSOvSNQ1SSGr2s0zfochfyh56tWJNmkcT1Pb4Qv6t5xOhZGm0V6hdAtg5
2wjfqXE4Rw44x+ycMEaYfFrxGxVAJgVKMIOqj8PeihPZBRm0dCT7wxqtEAufbmpbgH6EwQqlBrOA
ASkeBvGMBTvsODbPa+AgQGJep8V3TExUSVi2MHxtp5OGVKeU1JqA1jlQIZ7SC1tqOwIboLzUqPE9
oRKmT6gqsVYoEbTuvAr+xhXGoeY+LQF8SASlNW47zBiGeorjJICwCxp06fR2pLR8uWkkc3IP5PUd
4uTZhjy29I+KIR141389kU3RlY+14KEAYSZPJVDXFrjd0ue0rxM8x3KFJdBcx5t7Nep//HHMtm1V
f0m6ZNCyYFqYpmFM7BuXjApBovKHKzcLpFQB4LDEOIN8cVCKN/XB0UICt9/UoKkD3fN7M+WhLjbb
LrKb5UnKe3ZOklnPHbGdUmNK5lR4BO6pDlE+mwVJtO/bCfryap/5xNsKcGiJ8OSdZPJ5jUjfDbvS
PcxZgSp92VZg/lAeqOTiePA+Xejgt8YB2eJEAiloAv4gWYiwwYZ36jx24DFgLuIUp3O4lAQXfBGc
K0uMwwjWdHMCn8IifNG7iOIIwt1u8cCrgnpFLMOQT35WZcVY/+PX+TEAl0J4eRjN4+cqaXIeaDRW
9VztQyYxXilyRlL7mZyJsdkus2kPPy49Mz1RX5bHNiFaWcAtnk1VrKCKrKkqEJTEUTBQxVT7182C
Vyb9x1e8cnzNBanKQQnKTFunfSG6WFJOSGRRdb1T5Tle2os+z8gTqT+req1JA6ID++fDrKHMmvUn
f7v/RFVncQ+4C+AyKVn8V5//7y0GHc32pp34Rli4/FUOqLHXokJaKw+5AbuGAUTonejhoKAMT3M0
CuTDw3xS08NlNa6q4+Go9GnSohZGimIf43roA1bR1n3efcZG6qO8bsnKMMhg1jQj1x0bIb69wMs5
o799JZd3Lnj28OKJTPezy1QcFp7Wc11fT74SbB9npzc8O+LNJ0p5Ts2+ZOz1OJi+9dOu/5yknKkB
nvSaOJN2VmAK7orBR09x1FRfpG0BKgqneEaKOGOiU6XKMti4pjPr4yEguXycnyWzN7XUiTQ+hh9E
fMEQx5QA0tfhM4//s5zwqAsTvJM0XOpl9ut6cBn44hQz/ji4aAozzasgTlx0nUmTgAsahnhw+q8H
48tmTztwaPBI8L71ATg4TLJ41ZOz8/07IlVJHQ4v0v3y9cQ8qpEmipjrUET5pTkwk8kfZvuxyGM0
jiwkv2RNI5fa8rFzcuz9llfvcIv3HKWSS/zqowDw9WHWWr1ECnrZ3Ot/robgrN8FQVnlphtrLIYD
fCapH9Amg2Ld+roezOtSLHYkZIZOWpznj3/qNRDCcL1yNjWQjKG++SfAA2YMoCXMj8gwnMG70pTm
UYD6yqqi5OeiViA/T5C0T3IekmE60VpxHFbkIJmEm908dy/stVxMq7b0c1suySA7AgqTJy82rZZ2
9p1MASwYexo8x82favyZEirjTPrr/TQNgh5uMzTQVKnEOhFGwiS0vtsGfKEtXKzVq/GsTdCFL3aJ
2fUwbxmx+oyHX+x0nQpPYjdex3D7689pgqYCkGJLEgEIBINhvSNMZ092w02LucfGGMdUyjGxJpRw
cBAu15MaiRJiDwI6KOR4ddPhZ2tsbWiZ3G57wr2MGTtN1JGgubFAFtGgA61jwnIEXNPlQR73hV3W
mP0cc070VEKRyGuTct2Q1MrbaX2T2LhQxOLtmeOtmEWMPwiDYUdu++iS38z0eJ5SYZWTASAuSkuM
eSuiZ9DgGV3ohofBxOw1yR+EFl6u/DM/p2s5F+LkITJFiYu/jS+y28A76ylljpv/CeAITVJ5b/pu
pVx6bhOutRr+5mJAR6bxaNoFbe5WwTpWtEUBoK7FhCEpZynvyoFWxNVHgSIbUjqTX5oHRYK9PzBf
bBl/HLHy3QfFIg41UlemIgvhwCFCOZ0WzrpIXFD+cE191SK17CoEZ9xYJhrxXGumCI/0CdL2Sgnp
LLVQe9X9i0cyd6Xh+jk48jKaWC0qhaKo6u7blCPQa4Yxh4doS98mv92DZOl0KNBzpKml08ZsNOro
xfgKNBytR9t4r+buu2xVX5JubDZURSo7qD9LM8NoXclhkxnRpoFzRVJ8t+Jo1WNYQMLjdzFKInJ2
fkw9rhpWyQ3IP9OY6ebf9S3mf3ZvK4j9oq1gWZTqvGaGGUndxFta76VY+v6T/deG4KtnYk24luAI
uYS3XlD7e6N15VV0a8d59XRI00rZiEsetQ8jY5OUPHMWQZxYCVnHKnzuyTd9iu7fLJbp21Uwj/uV
wpF+tB3Z9kPPRPN9mYKuJoKwEiiF7guxvkDstUBcCh+arkxMmalTcV7YqJH7rhbORZPqULYNSD3B
HeZJFVvpWEQxBPL1xq9Z0vOdyk4sG1TdsU7jn3HhT9WjgywaT522j4xV/qfYLIvB7ig66on8iBXy
K+3ndvljL7hRmtyxjS5en6GRGBGXnRnQkCeMS0hpFTYMrngvVTUekHX4JxnBJi6JJgkBbO6mBDIt
El9uYMRuBp3ojt+hvomwdOczziiZTE9ALMoFzVanyiYt0Nb2Yi1EmqrqtMP7QvpvTV+T6tljgtC0
6PQzCxrCnZ/K530MexQeYgD12TqMWTG3wf727GIKguxHuXM8QhX7EV2FK4ZKVwE6SPK0tdpRFaWP
ZwaYfYvc7OYUiKsbzOMZVva8GOVdDAA955VwviDlDeMolSRzmwZwQQ4U/crXX81e57ybIawLNE0U
JZmBpMqtc5jBCZqtm1rlJq/7IMY8s9jAn/v1r9c5IAoa1ofkAvejWo07bm2PYUCTfdx3Y/0ajfy3
AgvHpD8oY2HmsKHmSBd10YfPL76QjEb8PCGgyvbFjHHiTszhZMBKhJOggmpHjannq+3PfB89yIT8
naykFbHkG22zuLOa+DgM0gyDRl920hbuA2mH46gzy7eQFVogmA475hPZmzIrMMlbGFiCHS7s2V64
TJEaVasAez0I6KUY1lamezYTCl/y8R+aczMU2Qo5Wadd9AN8sVG7hLH56QSdPdnbewGljnefVuGb
m9k8aQKqTapiz/c4CQk2p8P9HiaSbjsz/mlxUDm86IuGPKCrILwW2xs/GpNO6WvWuX5rw9GVRckL
Wv68SFPPJgh2uHHEPnrezQoVeC3S9NnqLT7W89ai/gbiZznY9uvB1VdKWiN24g36WXuU6pcr911B
IV+qQj4qT0IatFIukYJq4iq7c5PscauPCKnjH5TJYtMbpwBpMWntX6oXeRpXvhYLCcRd4YhwwXpC
XGdrxwAnj/5r2mq+6T+QxO9neQaYIArKm2WuUV0jDRdluYWxLaDWBPW8U2IlJxCE6fGY4RuHm/qT
bZpBsqcaaoW1C5GjKNTkZ2n94qsyBs6ZcZMdviTdiWsOYKr39WUzAZT6lEh1lorKSMmSdbEF3CoF
5S+BTh6DsSp0XZe+kR2mLVYrS+cv2UbkYuzNKxOAFNIy1+sHdwShSEkuF4sVbyOL2WqwkJW0Owq+
ZvLOTFAWDebLRMQpLadEmvfuibYHA600laBzEe4pWv1xGN6wnp1TVsL4iozdKF9OvrytNfJoF5Aj
lpoaTq8WekA+L3oEGHK2YSL/uKY9xOLKhs6lvUd8zx7F7SnnAG9iD2HONFvv7eeZtbG5koI9OdFP
V9gvzVGhHf9XMHFZAa5jeWkQ/IcrGO4v+rKC6LAetP8eYWICDnhDmhe2j2U+EGIk23uJtzhkClev
+EOWYBStufCFz1qID9UrB8gZL1O3XOBZaAwyXEZdVkEi3d7Zs0iW8noPgj59wR28Ht5/Revk4ovl
BgfZ1lHJ+i6M+4HTw5pIrBOCr+2GDTzpM8tNwhn5sZi3T7vuzBVEJEPLenOTcOaKPCETkgFoJDD7
d0gRX+jAUAVNfIHE227/1FHRUvUvq8PbtdFFcdCUM8u4ZAob8LC4sVXGexvbzX1wpMO9nZ5IsD/n
nTojIepXhaFemKp/51Tku++8363y8J6iPPt5Mjrwy524AYPjSeRh039eihNf4ZQdvcDO5q9Lwa/E
Aiun/MjVpaB2JqQxZfNeIPYTjCUBKDFcA0GmjSpqmc0MeD9zoerKZhvfGaXZQmgPeY0Fz8NiwWQo
R2KuXFs8mSKzIsENC+tG9Y1qt7Pg/032PzIuBveNm0GnjjOUizSDLcqJ+cXGrK6G84kBccg5RvdZ
aoX/g5yFu1IFMY9Vr+clivrh8wmFfkmDC6bQwayjFwt+76JAN1RIrKJyvVgPt5EmmOcQcwwXx4l2
hvQLNlXVXAg/AQjmB5SB3rBptvnUecTME4TDesoAi9efBYCuSKb3oJizM96E5xVhjSILcXTrxHjB
I7dVyqxXf3b7ZcZIaXfM0Kr0iSCYWRA4dW4Nxxt3huNiXB/6A5wbw6A8J1BIDrTOmEAOD9s8tZZE
MaCvR69vIIoCmXWRnskldOG000hL8uGuNmA030CYsX0zJWS+slY/VmLTFdPcjfZpswxcKwcObzl1
9YluA3n58PXErVIZepsr+a6i3SbSUWF/QSXpKpX2TZxdkFFZsiSBFFcvMpL+Yif6wQ1F6fTrduCA
aQLOhGcvJCSYWXaGQ6RQ4XCXYLFYFHZKYS/Q2WggMEdpBd8bVwK2osHNDSDW63AkWTvuRTlMSnUL
felWOddJz3QWE06a3OVBlr/i39nB0PXpy8bU5hGXKDG/NfxH9v57rGeEVDGwgwpq7nQhz9wyvcao
KVgrhIiNnDcPVoy6GXMBGMEvbg2xxLNWspmaUgrIQ3CDi9a6rhATveYB6T8kIsJlqRDpIfHdR30r
oD4NuAqtsIWqARwSBWpVxozhJp9JB1XaCDvHCcBT9rt210QlTptNH51DfYisonZzk13CJ75ZruoS
QAKWeQ7pVxux+/fR6DUQm3YIy93GK+zPXdXi42v/68pKCZ3GqmX+TcwqRvD2KWLi/FQQUjRzuSL2
L8/XwzVMuixe/PfhcUwKuso5ejA/8qil4ugIfvNWG0PG0dxg6BSfiF7LtiLFPSx7kjAz5ja3QGYE
Ap8m5gTpx8uP1hJCfQlEFaQv60PiXnJwBQbxQIQLix+pKvDAYUo9hqs9Yf9yoPA4QGgwq+hvwFEJ
L+S9k1aG6sPKOwAIZKh7VM2UDB9xdV5UvIBPGzJ+T2Wep+cCRU5mitfD/UnEmjLmFUc66pSoOVlY
zsRbVqjTIdhu7r+oFH8O4sL5VAVYanIqeazB4fMwg5qtw1otcsbXWcx/5uMhROdQQjHDP7jHRLjt
Cu9jMvdf05QisV0R1N4t5DP33bWvOOJScCnl/+CkVhxQWoHI5c8TI6wqMn2uwCoTynR5LZVDW9qe
Qwgib2p77YDvhEsKMBShFlacamWLaqxqq9GfrWegFgrUeNxaEQSdqMaVKxIxhpxIW0dhRsbCehFg
c10ly32wImPyCJQ3c+AwNNSBiZkhJZXJriTyddunIjigAuJsYqD1dpPd5BFYriw6Jg+Q2Y0B27Ou
sZo6ZD8igCP16bUTv3RzRz+/zqAbJ6uuUT/Ba3NEr9H/F/O6i4PI9bdKdGQwMyHmj3bR9rrNSBok
+ojrgqnLUpD2r9GMbHoFSN82GUDkf8QJJkX0k+mt1AceyCzddvC3dTxptBIrjb0rVmhyBA60iHSv
Dt7fy+GfCeOWYEKZpH6sFMTJcyApKG0z/zBvcOBze7WgAkdOUjDpwWEaBYiK/ibJn/PWZShOveiK
mvc4ee6NtH6EPzpLhFgc7YJnBXN4e0q4wjRUD/oSNo2cW1jnQ8Njmai4OpCDGJLKF2ebo8W3O9l+
s56/yZtReea7DxZDWE8Iej2Rctr3bpIF7hkTTetqpyffJJHer350SPkiDOqkUSnblW2W34+n0/wa
OHcVLYmfJJTuz9oSY8B4ploiUEMHvQMnzZ/jVIi9j2iXj8aQ/hngcqomi/4As0Yu8osSKPrWFlxn
reOVG4Ctxiovt7/ksODRqx/oXDXM3QXeEVGFAQdMKm2JtcX0RaANRxHZBTvrEkcagH6tWIgY6ksZ
1+t2M+84es8L+00o3fN8EY+8rr9H2avxFVoDde1TvpJhnRRgBS/5KSeubqvIQujEOc5FnP4o1cRT
r9b9Vqz2oR4ruO5Z9upwsUWRsB5VUxRbh5u6rwzGq3p7XpmQGYAVoxd419nZp9IesUf7sLjBbg2v
DoID7C6tGJzuuLhbTt4DaFp6qN2dgrc8fNP2UBeEaHF3p/98FspZq2v3gPYzyLiEOS7+NHs+qltT
O9GbxhKPxZ81QnfV/ytHasWyf0VPXHSrsblyOU7iPl7p5nDdWZc2FDk1Aigwn9nyqYn54xk2CXnO
L+UKSu+ixMy9poCaLV59+42Ab4fUjAPT+ZUUXwcXHhm3TGsQXhvjMUE4p1HHOOXKGmRFrIDPLqMS
kFFBiX6JprJWHrAHuarvDj05N19y2GHofOKHMaBfwYYomtovlyImM37ja6/RJmiwfyxxT+bJ+5NP
1Ecbo9bieDuBWC3HEfmCkHhY+dBxmVcgBdL6QvHonBQ8v8UoLzpw2uc5VlYRxkHPEWqGyEzAr8RS
Hsj076BiDvc4qOrzdNuRV7WmJarU8yYOQ4udIgLYmUFhAK2K1sCCY4Y7wkP+040TmjLPpmhGZxsk
KJmFUSuWhyKmHz3PQF1irKmd0HsHZZ9hQz4md+ELafu/MdLqfnJdUrhg0U/+pnB7xjRktsaT5s5+
VUDVHVOUvhJcNkN9gLVfCHe8Gn0tCXBOC/tXx6S4rQY/cFibsPkiyV1XcrJdXVmxc4xXWCrxDj3h
LG1xOrcwGVGOhaGRPD8ZPXQfuG4slKFMn6Vso4sbfHUSnd9LfHWyfkMeu/WEWylqT3s743J8p95l
HPPIGDztrWv/PmtNoszi+ssQ2bLZO/bjjhZ4CpKoxfDxLiYFTDrqh5eag+SXA9uJl2qytldYmXus
zMffEZDEHnpas9ldtVKL2zUQTA1hjNg+dT87Ho0F1ld0Q9UnOtGVx0Hjvdv0ySqHsgRCclyd7kWD
DNDqU21GRcuVFacYFoE9wjWExSjMTBS3JCLpVe87yweZ2Uvt8ORsM7fhRbLMT84T1861NUNIWd41
Cs211vufkXbhVX2GbRv7kfDvI6iedZZym7qE/yleHJgyz40EpTiHez9jMqwJOcjCt31wh1AJGIXp
DpASyklb5//t253NVP9gIKRJN7is4GkAc+XshjRz/ieSko9nJb0Uy3oND60W46xA8lg4ife4zAwG
nfk2h2MUS3LGmgqHEk6LqbUk/tg1BUO2t3Zc9zjJjosYdJ+IIaw9sH02Fn87oY6hE+scGN8axPag
teAIvAugHmRe2zoNXbnVEtUGAxtPwHteOxf1J0opxylB8CbMuK2LrPTNTe544jAcxUC3M/OcbFEq
A5Lj6haomHeNvEJhnxjdvYQSMQk+WyPNH0Btg3+NjKSsC8QesqO9S0LSjoBf4UimFbvnsgZ5+bRU
/OY5SGmPkyy4fWlCT9U1qXHK0aF/porhHZUtX9qoOOYhQH9oaASpp6mKr5wnx5t/ZaUmeOTLXQX9
9k5XwlRlCr+rbAxR9q7ukCf+pnHVSOLhTfMEEerpowhWp74YRt3xqoEuAX2XE9/PAKkP23rTNDXW
bWQSwkpL/AKYKx66uhTXiVVVD9EvLgfsMZxcOInSDBCt/rkap2rMLTfAZxdcMwfFlujyRj92GaZ2
unRbVQidzMXdQEc2XC+R3Iv+nBOIu7S5WnfNme1x6IarQfUlpUEPcCLUC2juGsHyGsf50+2ef8pc
wNLVMOjZ1+zgzd++K79HbAeBGD4Z8iZPfAP7QMRJPVhY3jHQ9zMiDt0d2MSjjt94BwisjDIY2gHd
+SqhTNmMqEdPDNwAu0gBO020kr7Z76W/834lZ0yTXHEzh2ujAwlu93a9UeaaH0PxNgCfZoqI6rEm
EoDUkafpEIGi7zSdW0GCI3yZapyDhn6jQc24vTC2qLMU96BTKjzwqAczNshpn2ZJC+kjTbh0b4L9
uFqrtjIaEylw6ImKFh3gQoHDd2bH6slsF/Cu2p5cSj6dAzaetEk43E76xV3FNWh8mek5x6SpGXdd
eobISHttNr9BT655Zcpyx2qYl9BivjutmeeMAOl3f8rogaUuAQh3XsPhPMaoK3MCaHQHDZA5dOC1
QA67FQ4krVAJ7XjDSd3pIDoQTaHX+gNHEK7R8ZthM8VOBuilbhMl6LVqzFSNVSJQB5JDnU9AFe4b
vcYIGuuto38hBGpBAEnsXJXoiDdeOzoSK8mvCSr+2ut/1WJsA4MLuUGRPIYRZyBAkhi4rdimqBRl
wB+z5ZgYlvGBofV63/vz87HLWk2Lz8CmAQFBwq1p0kQhoNns5wxe/S5HJ+1UCB1x6t3LyFSPebPh
-- ==============================================================
-- RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
-- Version: 2020.1
-- Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
-- 
-- ===========================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity myproject is
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    fc1_input_V_ap_vld : IN STD_LOGIC;
    fc1_input_V : IN STD_LOGIC_VECTOR (255 downto 0);
    layer13_out_0_V : OUT STD_LOGIC_VECTOR (15 downto 0);
    layer13_out_0_V_ap_vld : OUT STD_LOGIC;
    layer13_out_1_V : OUT STD_LOGIC_VECTOR (15 downto 0);
    layer13_out_1_V_ap_vld : OUT STD_LOGIC;
    layer13_out_2_V : OUT STD_LOGIC_VECTOR (15 downto 0);
    layer13_out_2_V_ap_vld : OUT STD_LOGIC;
    layer13_out_3_V : OUT STD_LOGIC_VECTOR (15 downto 0);
    layer13_out_3_V_ap_vld : OUT STD_LOGIC;
    layer13_out_4_V : OUT STD_LOGIC_VECTOR (15 downto 0);
    layer13_out_4_V_ap_vld : OUT STD_LOGIC;
    const_size_in_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
    const_size_in_1_ap_vld : OUT STD_LOGIC;
    const_size_out_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
    const_size_out_1_ap_vld : OUT STD_LOGIC );
end;


architecture behav of myproject is 
    attribute CORE_GENERATION_INFO : STRING;
    attribute CORE_GENERATION_INFO of behav : architecture is
    "myproject,hls_ip_2020_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7vx415t-ffg1157-1,HLS_INPUT_CLOCK=5.000000,HLS_INPUT_ARCH=pipeline,HLS_SYN_CLOCK=4.367250,HLS_SYN_LAT=38,HLS_SYN_TPT=1,HLS_SYN_MEM=4,HLS_SYN_DSP=2808,HLS_SYN_FF=272473,HLS_SYN_LUT=113927,HLS_VERSION=2020_1}";
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';
    constant ap_ST_fsm_pp0_stage0 : STD_LOGIC_VECTOR (0 downto 0) := "1";
    constant ap_const_lv32_0 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000000";
    constant ap_const_boolean_1 : BOOLEAN := true;
    constant ap_const_boolean_0 : BOOLEAN := false;
    constant ap_const_lv256_lc_1 : STD_LOGIC_VECTOR (255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_const_lv16_10 : STD_LOGIC_VECTOR (15 downto 0) := "0000000000010000";
    constant ap_const_lv16_5 : STD_LOGIC_VECTOR (15 downto 0) := "0000000000000101";

    signal ap_CS_fsm : STD_LOGIC_VECTOR (0 downto 0) := "1";
    attribute fsm_encoding : string;
    attribute fsm_encoding of ap_CS_fsm : signal is "none";
    signal ap_CS_fsm_pp0_stage0 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage0 : signal is "none";
    signal ap_enable_reg_pp0_iter0 : STD_LOGIC;
    signal ap_enable_reg_pp0_iter1 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter2 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter3 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter4 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter5 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter6 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter7 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter8 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter9 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter10 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter11 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter12 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter13 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter14 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter15 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter16 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter17 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter18 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter19 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter20 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter21 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter22 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter23 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter24 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter25 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter26 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter27 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter28 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter29 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter30 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter31 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter32 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter33 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter34 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter35 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter36 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter37 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter38 : STD_LOGIC := '0';
    signal ap_idle_pp0 : STD_LOGIC;
    signal fc1_input_V_ap_vld_in_sig : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10 : BOOLEAN;
    signal ap_block_state12_pp0_stage0_iter11 : BOOLEAN;
    signal ap_block_state13_pp0_stage0_iter12 : BOOLEAN;
    signal ap_block_state14_pp0_stage0_iter13 : BOOLEAN;
    signal ap_block_state15_pp0_stage0_iter14 : BOOLEAN;
    signal ap_block_state16_pp0_stage0_iter15 : BOOLEAN;
    signal ap_block_state17_pp0_stage0_iter16 : BOOLEAN;
    signal ap_block_state18_pp0_stage0_iter17 : BOOLEAN;
    signal ap_block_state19_pp0_stage0_iter18 : BOOLEAN;
    signal ap_block_state20_pp0_stage0_iter19 : BOOLEAN;
    signal ap_block_state21_pp0_stage0_iter20 : BOOLEAN;
    signal ap_block_state22_pp0_stage0_iter21 : BOOLEAN;
    signal ap_block_state23_pp0_stage0_iter22 : BOOLEAN;
    signal ap_block_state24_pp0_stage0_iter23 : BOOLEAN;
    signal ap_block_state25_pp0_stage0_iter24 : BOOLEAN;
    signal ap_block_state26_pp0_stage0_iter25 : BOOLEAN;
    signal ap_block_state27_pp0_stage0_iter26 : BOOLEAN;
    signal ap_block_state28_pp0_stage0_iter27 : BOOLEAN;
    signal ap_block_state29_pp0_stage0_iter28 : BOOLEAN;
    signal ap_block_state30_pp0_stage0_iter29 : BOOLEAN;
    signal ap_block_state31_pp0_stage0_iter30 : BOOLEAN;
    signal ap_block_state32_pp0_stage0_iter31 : BOOLEAN;
    signal ap_block_state33_pp0_stage0_iter32 : BOOLEAN;
    signal ap_block_state34_pp0_stage0_iter33 : BOOLEAN;
    signal ap_block_state35_pp0_stage0_iter34 : BOOLEAN;
    signal ap_block_state36_pp0_stage0_iter35 : BOOLEAN;
    signal ap_block_state37_pp0_stage0_iter36 : BOOLEAN;
    signal ap_block_state38_pp0_stage0_iter37 : BOOLEAN;
    signal ap_block_state39_pp0_stage0_iter38 : BOOLEAN;
    signal ap_block_pp0_stage0_11001 : BOOLEAN;
    signal fc1_input_V_preg : STD_LOGIC_VECTOR (255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    signal fc1_input_V_in_sig : STD_LOGIC_VECTOR (255 downto 0);
    signal fc1_input_V_ap_vld_preg : STD_LOGIC := '0';
    signal fc1_input_V_blk_n : STD_LOGIC;
    signal ap_block_pp0_stage0 : BOOLEAN;
    signal layer2_out_0_V_reg_1501 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_1_V_reg_1506 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_2_V_reg_1511 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_3_V_reg_1516 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_4_V_reg_1521 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_5_V_reg_1526 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_6_V_reg_1531 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_7_V_reg_1536 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_8_V_reg_1541 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_9_V_reg_1546 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_10_V_reg_1551 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_11_V_reg_1556 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_12_V_reg_1561 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_13_V_reg_1566 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_14_V_reg_1571 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_15_V_reg_1576 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_16_V_reg_1581 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_17_V_reg_1586 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_18_V_reg_1591 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_19_V_reg_1596 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_20_V_reg_1601 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_21_V_reg_1606 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_22_V_reg_1611 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_23_V_reg_1616 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_24_V_reg_1621 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_25_V_reg_1626 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_26_V_reg_1631 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_27_V_reg_1636 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_28_V_reg_1641 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_29_V_reg_1646 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_30_V_reg_1651 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_31_V_reg_1656 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_32_V_reg_1661 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_33_V_reg_1666 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_34_V_reg_1671 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_35_V_reg_1676 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_36_V_reg_1681 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_37_V_reg_1686 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_38_V_reg_1691 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_39_V_reg_1696 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_40_V_reg_1701 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_41_V_reg_1706 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_42_V_reg_1711 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_43_V_reg_1716 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_44_V_reg_1721 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_45_V_reg_1726 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_46_V_reg_1731 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_47_V_reg_1736 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_48_V_reg_1741 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_49_V_reg_1746 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_50_V_reg_1751 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_51_V_reg_1756 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_52_V_reg_1761 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_53_V_reg_1766 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_54_V_reg_1771 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_55_V_reg_1776 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_56_V_reg_1781 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_57_V_reg_1786 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_58_V_reg_1791 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_59_V_reg_1796 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_60_V_reg_1801 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_61_V_reg_1806 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_62_V_reg_1811 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer2_out_63_V_reg_1816 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_0_V_reg_1821 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_1_V_reg_1826 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_2_V_reg_1831 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_3_V_reg_1836 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_4_V_reg_1841 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_5_V_reg_1846 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_6_V_reg_1851 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_7_V_reg_1856 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_8_V_reg_1861 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_9_V_reg_1866 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_10_V_reg_1871 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_11_V_reg_1876 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_12_V_reg_1881 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_13_V_reg_1886 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_14_V_reg_1891 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_15_V_reg_1896 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_16_V_reg_1901 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_17_V_reg_1906 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_18_V_reg_1911 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_19_V_reg_1916 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_20_V_reg_1921 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_21_V_reg_1926 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_22_V_reg_1931 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_23_V_reg_1936 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_24_V_reg_1941 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_25_V_reg_1946 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_26_V_reg_1951 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_27_V_reg_1956 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_28_V_reg_1961 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_29_V_reg_1966 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_30_V_reg_1971 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_31_V_reg_1976 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_32_V_reg_1981 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_33_V_reg_1986 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_34_V_reg_1991 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_35_V_reg_1996 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_36_V_reg_2001 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_37_V_reg_2006 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_38_V_reg_2011 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_39_V_reg_2016 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_40_V_reg_2021 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_41_V_reg_2026 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_42_V_reg_2031 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_43_V_reg_2036 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_44_V_reg_2041 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_45_V_reg_2046 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_46_V_reg_2051 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_47_V_reg_2056 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_48_V_reg_2061 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_49_V_reg_2066 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_50_V_reg_2071 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_51_V_reg_2076 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_52_V_reg_2081 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_53_V_reg_2086 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_54_V_reg_2091 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_55_V_reg_2096 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_56_V_reg_2101 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_57_V_reg_2106 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_58_V_reg_2111 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_59_V_reg_2116 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_60_V_reg_2121 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_61_V_reg_2126 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_62_V_reg_2131 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer4_out_63_V_reg_2136 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_0_V_reg_2141 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_1_V_reg_2146 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_2_V_reg_2151 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_3_V_reg_2156 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_4_V_reg_2161 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_5_V_reg_2166 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_6_V_reg_2171 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_7_V_reg_2176 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_8_V_reg_2181 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_9_V_reg_2186 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_10_V_reg_2191 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_11_V_reg_2196 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_12_V_reg_2201 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_13_V_reg_2206 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_14_V_reg_2211 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_15_V_reg_2216 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_16_V_reg_2221 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_17_V_reg_2226 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_18_V_reg_2231 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_19_V_reg_2236 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_20_V_reg_2241 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_21_V_reg_2246 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_22_V_reg_2251 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_23_V_reg_2256 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_24_V_reg_2261 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_25_V_reg_2266 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_26_V_reg_2271 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_27_V_reg_2276 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_28_V_reg_2281 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_29_V_reg_2286 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_30_V_reg_2291 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer5_out_31_V_reg_2296 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_0_V_reg_2301 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_1_V_reg_2306 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_2_V_reg_2311 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_3_V_reg_2316 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_4_V_reg_2321 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_5_V_reg_2326 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_6_V_reg_2331 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_7_V_reg_2336 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_8_V_reg_2341 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_9_V_reg_2346 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_10_V_reg_2351 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_11_V_reg_2356 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_12_V_reg_2361 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_13_V_reg_2366 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_14_V_reg_2371 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_15_V_reg_2376 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_16_V_reg_2381 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_17_V_reg_2386 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_18_V_reg_2391 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_19_V_reg_2396 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_20_V_reg_2401 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_21_V_reg_2406 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_22_V_reg_2411 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_23_V_reg_2416 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_24_V_reg_2421 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_25_V_reg_2426 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_26_V_reg_2431 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_27_V_reg_2436 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_28_V_reg_2441 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_29_V_reg_2446 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_30_V_reg_2451 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer7_out_31_V_reg_2456 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_0_V_reg_2461 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_1_V_reg_2466 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_2_V_reg_2471 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_3_V_reg_2476 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_4_V_reg_2481 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_5_V_reg_2486 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_6_V_reg_2491 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_7_V_reg_2496 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_8_V_reg_2501 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_9_V_reg_2506 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_10_V_reg_2511 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_11_V_reg_2516 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_12_V_reg_2521 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_13_V_reg_2526 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_14_V_reg_2531 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_15_V_reg_2536 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_16_V_reg_2541 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_17_V_reg_2546 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_18_V_reg_2551 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_19_V_reg_2556 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_20_V_reg_2561 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_21_V_reg_2566 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_22_V_reg_2571 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_23_V_reg_2576 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_24_V_reg_2581 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_25_V_reg_2586 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_26_V_reg_2591 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_27_V_reg_2596 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_28_V_reg_2601 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_29_V_reg_2606 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_30_V_reg_2611 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer8_out_31_V_reg_2616 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_0_V_reg_2621 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_1_V_reg_2626 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_2_V_reg_2631 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_3_V_reg_2636 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_4_V_reg_2641 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_5_V_reg_2646 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_6_V_reg_2651 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_7_V_reg_2656 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_8_V_reg_2661 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_9_V_reg_2666 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_10_V_reg_2671 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_11_V_reg_2676 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_12_V_reg_2681 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_13_V_reg_2686 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_14_V_reg_2691 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_15_V_reg_2696 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_16_V_reg_2701 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_17_V_reg_2706 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_18_V_reg_2711 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_19_V_reg_2716 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_20_V_reg_2721 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_21_V_reg_2726 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_22_V_reg_2731 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_23_V_reg_2736 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_24_V_reg_2741 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_25_V_reg_2746 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_26_V_reg_2751 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_27_V_reg_2756 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_28_V_reg_2761 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_29_V_reg_2766 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_30_V_reg_2771 : STD_LOGIC_VECTOR (15 downto 0);
    signal layer10_out_31_V_reg_2776 : STD_LOGIC_VECTOR (15 downto 0);
    signal ap_block_pp0_stage0_subdone : BOOLEAN;
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call145 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call145 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call145 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call145 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call145 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call145 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call145 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call145 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call145 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9_ignore_call145 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10_ignore_call145 : BOOLEAN;
    signal ap_block_state12_pp0_stage0_iter11_ignore_call145 : BOOLEAN;
    signal ap_block_state13_pp0_stage0_iter12_ignore_call145 : BOOLEAN;
    signal ap_block_state14_pp0_stage0_iter13_ignore_call145 : BOOLEAN;
    signal ap_block_state15_pp0_stage0_iter14_ignore_call145 : BOOLEAN;
    signal ap_block_state16_pp0_stage0_iter15_ignore_call145 : BOOLEAN;
    signal ap_block_state17_pp0_stage0_iter16_ignore_call145 : BOOLEAN;
    signal ap_block_state18_pp0_stage0_iter17_ignore_call145 : BOOLEAN;
    signal ap_block_state19_pp0_stage0_iter18_ignore_call145 : BOOLEAN;
    signal ap_block_state20_pp0_stage0_iter19_ignore_call145 : BOOLEAN;
    signal ap_block_state21_pp0_stage0_iter20_ignore_call145 : BOOLEAN;
    signal ap_block_state22_pp0_stage0_iter21_ignore_call145 : BOOLEAN;
    signal ap_block_state23_pp0_stage0_iter22_ignore_call145 : BOOLEAN;
    signal ap_block_state24_pp0_stage0_iter23_ignore_call145 : BOOLEAN;
    signal ap_block_state25_pp0_stage0_iter24_ignore_call145 : BOOLEAN;
    signal ap_block_state26_pp0_stage0_iter25_ignore_call145 : BOOLEAN;
    signal ap_block_state27_pp0_stage0_iter26_ignore_call145 : BOOLEAN;
    signal ap_block_state28_pp0_stage0_iter27_ignore_call145 : BOOLEAN;
    signal ap_block_state29_pp0_stage0_iter28_ignore_call145 : BOOLEAN;
    signal ap_block_state30_pp0_stage0_iter29_ignore_call145 : BOOLEAN;
    signal ap_block_state31_pp0_stage0_iter30_ignore_call145 : BOOLEAN;
    signal ap_block_state32_pp0_stage0_iter31_ignore_call145 : BOOLEAN;
    signal ap_block_state33_pp0_stage0_iter32_ignore_call145 : BOOLEAN;
    signal ap_block_state34_pp0_stage0_iter33_ignore_call145 : BOOLEAN;
    signal ap_block_state35_pp0_stage0_iter34_ignore_call145 : BOOLEAN;
    signal ap_block_state36_pp0_stage0_iter35_ignore_call145 : BOOLEAN;
    signal ap_block_state37_pp0_stage0_iter36_ignore_call145 : BOOLEAN;
    signal ap_block_state38_pp0_stage0_iter37_ignore_call145 : BOOLEAN;
    signal ap_block_state39_pp0_stage0_iter38_ignore_call145 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp177 : BOOLEAN;
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_32 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_33 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_34 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_35 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_36 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_37 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_38 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_39 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_40 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_41 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_42 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_43 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_44 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_45 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_46 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_47 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_48 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_49 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_50 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_51 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_52 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_53 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_54 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_55 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_56 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_57 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_58 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_59 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_60 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_61 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_62 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_63 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call15 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call15 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call15 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call15 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call15 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call15 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call15 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call15 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call15 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9_ignore_call15 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10_ignore_call15 : BOOLEAN;
    signal ap_block_state12_pp0_stage0_iter11_ignore_call15 : BOOLEAN;
    signal ap_block_state13_pp0_stage0_iter12_ignore_call15 : BOOLEAN;
    signal ap_block_state14_pp0_stage0_iter13_ignore_call15 : BOOLEAN;
    signal ap_block_state15_pp0_stage0_iter14_ignore_call15 : BOOLEAN;
    signal ap_block_state16_pp0_stage0_iter15_ignore_call15 : BOOLEAN;
    signal ap_block_state17_pp0_stage0_iter16_ignore_call15 : BOOLEAN;
    signal ap_block_state18_pp0_stage0_iter17_ignore_call15 : BOOLEAN;
    signal ap_block_state19_pp0_stage0_iter18_ignore_call15 : BOOLEAN;
    signal ap_block_state20_pp0_stage0_iter19_ignore_call15 : BOOLEAN;
    signal ap_block_state21_pp0_stage0_iter20_ignore_call15 : BOOLEAN;
    signal ap_block_state22_pp0_stage0_iter21_ignore_call15 : BOOLEAN;
    signal ap_block_state23_pp0_stage0_iter22_ignore_call15 : BOOLEAN;
    signal ap_block_state24_pp0_stage0_iter23_ignore_call15 : BOOLEAN;
    signal ap_block_state25_pp0_stage0_iter24_ignore_call15 : BOOLEAN;
    signal ap_block_state26_pp0_stage0_iter25_ignore_call15 : BOOLEAN;
    signal ap_block_state27_pp0_stage0_iter26_ignore_call15 : BOOLEAN;
    signal ap_block_state28_pp0_stage0_iter27_ignore_call15 : BOOLEAN;
    signal ap_block_state29_pp0_stage0_iter28_ignore_call15 : BOOLEAN;
    signal ap_block_state30_pp0_stage0_iter29_ignore_call15 : BOOLEAN;
    signal ap_block_state31_pp0_stage0_iter30_ignore_call15 : BOOLEAN;
    signal ap_block_state32_pp0_stage0_iter31_ignore_call15 : BOOLEAN;
    signal ap_block_state33_pp0_stage0_iter32_ignore_call15 : BOOLEAN;
    signal ap_block_state34_pp0_stage0_iter33_ignore_call15 : BOOLEAN;
    signal ap_block_state35_pp0_stage0_iter34_ignore_call15 : BOOLEAN;
    signal ap_block_state36_pp0_stage0_iter35_ignore_call15 : BOOLEAN;
    signal ap_block_state37_pp0_stage0_iter36_ignore_call15 : BOOLEAN;
    signal ap_block_state38_pp0_stage0_iter37_ignore_call15 : BOOLEAN;
    signal ap_block_state39_pp0_stage0_iter38_ignore_call15 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp41 : BOOLEAN;
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call211 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call211 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call211 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call211 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call211 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call211 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call211 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call211 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call211 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9_ignore_call211 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10_ignore_call211 : BOOLEAN;
    signal ap_block_state12_pp0_stage0_iter11_ignore_call211 : BOOLEAN;
    signal ap_block_state13_pp0_stage0_iter12_ignore_call211 : BOOLEAN;
    signal ap_block_state14_pp0_stage0_iter13_ignore_call211 : BOOLEAN;
    signal ap_block_state15_pp0_stage0_iter14_ignore_call211 : BOOLEAN;
    signal ap_block_state16_pp0_stage0_iter15_ignore_call211 : BOOLEAN;
    signal ap_block_state17_pp0_stage0_iter16_ignore_call211 : BOOLEAN;
    signal ap_block_state18_pp0_stage0_iter17_ignore_call211 : BOOLEAN;
    signal ap_block_state19_pp0_stage0_iter18_ignore_call211 : BOOLEAN;
    signal ap_block_state20_pp0_stage0_iter19_ignore_call211 : BOOLEAN;
    signal ap_block_state21_pp0_stage0_iter20_ignore_call211 : BOOLEAN;
    signal ap_block_state22_pp0_stage0_iter21_ignore_call211 : BOOLEAN;
    signal ap_block_state23_pp0_stage0_iter22_ignore_call211 : BOOLEAN;
    signal ap_block_state24_pp0_stage0_iter23_ignore_call211 : BOOLEAN;
    signal ap_block_state25_pp0_stage0_iter24_ignore_call211 : BOOLEAN;
    signal ap_block_state26_pp0_stage0_iter25_ignore_call211 : BOOLEAN;
    signal ap_block_state27_pp0_stage0_iter26_ignore_call211 : BOOLEAN;
    signal ap_block_state28_pp0_stage0_iter27_ignore_call211 : BOOLEAN;
    signal ap_block_state29_pp0_stage0_iter28_ignore_call211 : BOOLEAN;
    signal ap_block_state30_pp0_stage0_iter29_ignore_call211 : BOOLEAN;
    signal ap_block_state31_pp0_stage0_iter30_ignore_call211 : BOOLEAN;
    signal ap_block_state32_pp0_stage0_iter31_ignore_call211 : BOOLEAN;
    signal ap_block_state33_pp0_stage0_iter32_ignore_call211 : BOOLEAN;
    signal ap_block_state34_pp0_stage0_iter33_ignore_call211 : BOOLEAN;
    signal ap_block_state35_pp0_stage0_iter34_ignore_call211 : BOOLEAN;
    signal ap_block_state36_pp0_stage0_iter35_ignore_call211 : BOOLEAN;
    signal ap_block_state37_pp0_stage0_iter36_ignore_call211 : BOOLEAN;
    signal ap_block_state38_pp0_stage0_iter37_ignore_call211 : BOOLEAN;
    signal ap_block_state39_pp0_stage0_iter38_ignore_call211 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp250 : BOOLEAN;
    signal grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_ce : STD_LOGIC;
    signal ap_block_state1_pp0_stage0_iter0_ignore_call277 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call277 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call277 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call277 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call277 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call277 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call277 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call277 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call277 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9_ignore_call277 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10_ignore_call277 : BOOLEAN;
    signal ap_block_state12_pp0_stage0_iter11_ignore_call277 : BOOLEAN;
    signal ap_block_state13_pp0_stage0_iter12_ignore_call277 : BOOLEAN;
    signal ap_block_state14_pp0_stage0_iter13_ignore_call277 : BOOLEAN;
    signal ap_block_state15_pp0_stage0_iter14_ignore_call277 : BOOLEAN;
    signal ap_block_state16_pp0_stage0_iter15_ignore_call277 : BOOLEAN;
    signal ap_block_state17_pp0_stage0_iter16_ignore_call277 : BOOLEAN;
    signal ap_block_state18_pp0_stage0_iter17_ignore_call277 : BOOLEAN;
    signal ap_block_state19_pp0_stage0_iter18_ignore_call277 : BOOLEAN;
    signal ap_block_state20_pp0_stage0_iter19_ignore_call277 : BOOLEAN;
    signal ap_block_state21_pp0_stage0_iter20_ignore_call277 : BOOLEAN;
    signal ap_block_state22_pp0_stage0_iter21_ignore_call277 : BOOLEAN;
    signal ap_block_state23_pp0_stage0_iter22_ignore_call277 : BOOLEAN;
    signal ap_block_state24_pp0_stage0_iter23_ignore_call277 : BOOLEAN;
    signal ap_block_state25_pp0_stage0_iter24_ignore_call277 : BOOLEAN;
    signal ap_block_state26_pp0_stage0_iter25_ignore_call277 : BOOLEAN;
    signal ap_block_state27_pp0_stage0_iter26_ignore_call277 : BOOLEAN;
    signal ap_block_state28_pp0_stage0_iter27_ignore_call277 : BOOLEAN;
    signal ap_block_state29_pp0_stage0_iter28_ignore_call277 : BOOLEAN;
    signal ap_block_state30_pp0_stage0_iter29_ignore_call277 : BOOLEAN;
    signal ap_block_state31_pp0_stage0_iter30_ignore_call277 : BOOLEAN;
    signal ap_block_state32_pp0_stage0_iter31_ignore_call277 : BOOLEAN;
    signal ap_block_state33_pp0_stage0_iter32_ignore_call277 : BOOLEAN;
    signal ap_block_state34_pp0_stage0_iter33_ignore_call277 : BOOLEAN;
    signal ap_block_state35_pp0_stage0_iter34_ignore_call277 : BOOLEAN;
    signal ap_block_state36_pp0_stage0_iter35_ignore_call277 : BOOLEAN;
    signal ap_block_state37_pp0_stage0_iter36_ignore_call277 : BOOLEAN;
    signal ap_block_state38_pp0_stage0_iter37_ignore_call277 : BOOLEAN;
    signal ap_block_state39_pp0_stage0_iter38_ignore_call277 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp322 : BOOLEAN;
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_ready : STD_LOGIC;
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_32 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_33 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_34 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_35 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_36 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_37 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_38 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_39 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_40 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_41 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_42 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_43 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_44 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_45 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_46 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_47 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_48 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_49 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_50 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_51 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_52 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_53 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_54 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_55 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_56 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_57 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_58 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_59 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_60 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_61 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_62 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_63 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_ready : STD_LOGIC;
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_ready : STD_LOGIC;
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_5 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_6 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_7 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_8 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_9 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_10 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_11 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_12 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_13 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_14 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_15 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_16 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_17 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_18 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_19 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_20 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_21 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_22 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_23 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_24 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_25 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_26 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_27 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_28 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_29 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_30 : STD_LOGIC_VECTOR (15 downto 0);
    signal call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_31 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_done : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_idle : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_ready : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_ce : STD_LOGIC;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_1 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_2 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_3 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_4 : STD_LOGIC_VECTOR (15 downto 0);
    signal ap_block_state1_pp0_stage0_iter0_ignore_call283 : BOOLEAN;
    signal ap_block_state2_pp0_stage0_iter1_ignore_call283 : BOOLEAN;
    signal ap_block_state3_pp0_stage0_iter2_ignore_call283 : BOOLEAN;
    signal ap_block_state4_pp0_stage0_iter3_ignore_call283 : BOOLEAN;
    signal ap_block_state5_pp0_stage0_iter4_ignore_call283 : BOOLEAN;
    signal ap_block_state6_pp0_stage0_iter5_ignore_call283 : BOOLEAN;
    signal ap_block_state7_pp0_stage0_iter6_ignore_call283 : BOOLEAN;
    signal ap_block_state8_pp0_stage0_iter7_ignore_call283 : BOOLEAN;
    signal ap_block_state9_pp0_stage0_iter8_ignore_call283 : BOOLEAN;
    signal ap_block_state10_pp0_stage0_iter9_ignore_call283 : BOOLEAN;
    signal ap_block_state11_pp0_stage0_iter10_ignore_call283 : BOOLEAN;
    signal ap_block_state12_pp0_stage0_iter11_ignore_call283 : BOOLEAN;
    signal ap_block_state13_pp0_stage0_iter12_ignore_call283 : BOOLEAN;
    signal ap_block_state14_pp0_stage0_iter13_ignore_call283 : BOOLEAN;
    signal ap_block_state15_pp0_stage0_iter14_ignore_call283 : BOOLEAN;
    signal ap_block_state16_pp0_stage0_iter15_ignore_call283 : BOOLEAN;
    signal ap_block_state17_pp0_stage0_iter16_ignore_call283 : BOOLEAN;
    signal ap_block_state18_pp0_stage0_iter17_ignore_call283 : BOOLEAN;
    signal ap_block_state19_pp0_stage0_iter18_ignore_call283 : BOOLEAN;
    signal ap_block_state20_pp0_stage0_iter19_ignore_call283 : BOOLEAN;
    signal ap_block_state21_pp0_stage0_iter20_ignore_call283 : BOOLEAN;
    signal ap_block_state22_pp0_stage0_iter21_ignore_call283 : BOOLEAN;
    signal ap_block_state23_pp0_stage0_iter22_ignore_call283 : BOOLEAN;
    signal ap_block_state24_pp0_stage0_iter23_ignore_call283 : BOOLEAN;
    signal ap_block_state25_pp0_stage0_iter24_ignore_call283 : BOOLEAN;
    signal ap_block_state26_pp0_stage0_iter25_ignore_call283 : BOOLEAN;
    signal ap_block_state27_pp0_stage0_iter26_ignore_call283 : BOOLEAN;
    signal ap_block_state28_pp0_stage0_iter27_ignore_call283 : BOOLEAN;
    signal ap_block_state29_pp0_stage0_iter28_ignore_call283 : BOOLEAN;
    signal ap_block_state30_pp0_stage0_iter29_ignore_call283 : BOOLEAN;
    signal ap_block_state31_pp0_stage0_iter30_ignore_call283 : BOOLEAN;
    signal ap_block_state32_pp0_stage0_iter31_ignore_call283 : BOOLEAN;
    signal ap_block_state33_pp0_stage0_iter32_ignore_call283 : BOOLEAN;
    signal ap_block_state34_pp0_stage0_iter33_ignore_call283 : BOOLEAN;
    signal ap_block_state35_pp0_stage0_iter34_ignore_call283 : BOOLEAN;
    signal ap_block_state36_pp0_stage0_iter35_ignore_call283 : BOOLEAN;
    signal ap_block_state37_pp0_stage0_iter36_ignore_call283 : BOOLEAN;
    signal ap_block_state38_pp0_stage0_iter37_ignore_call283 : BOOLEAN;
    signal ap_block_state39_pp0_stage0_iter38_ignore_call283 : BOOLEAN;
    signal ap_block_pp0_stage0_11001_ignoreCallOp334 : BOOLEAN;
    signal grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start_reg : STD_LOGIC := '0';
    signal ap_block_pp0_stage0_01001 : BOOLEAN;
    signal ap_NS_fsm : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_idle_pp0_0to37 : STD_LOGIC;
    signal ap_reset_idle_pp0 : STD_LOGIC;
    signal ap_enable_pp0 : STD_LOGIC;

    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_32_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_33_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_34_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_35_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_36_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_37_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_38_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_39_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_40_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_41_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_42_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_43_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_44_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_45_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_46_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_47_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_48_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_49_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_50_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_51_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_52_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_53_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_54_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_55_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_56_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_57_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_58_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_59_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_60_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_61_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_62_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_63_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2 IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_V_read : IN STD_LOGIC_VECTOR (255 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_32 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_33 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_34 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_35 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_36 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_37 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_38 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_39 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_40 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_41 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_42 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_43 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_44 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_45 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_46 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_47 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_48 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_49 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_50 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_51 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_52 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_53 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_54 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_55 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_56 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_57 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_58 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_59 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_60 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_61 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_62 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_63 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0 IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_ce : IN STD_LOGIC );
    end component;


    component relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_32_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_33_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_34_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_35_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_36_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_37_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_38_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_39_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_40_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_41_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_42_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_43_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_44_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_45_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_46_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_47_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_48_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_49_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_50_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_51_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_52_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_53_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_54_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_55_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_56_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_57_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_58_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_59_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_60_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_61_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_62_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_63_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_32 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_33 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_34 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_35 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_36 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_37 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_38 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_39 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_40 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_41 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_42 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_43 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_44 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_45 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_46 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_47 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_48 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_49 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_50 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_51 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_52 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_53 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_54 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_55 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_56 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_57 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_58 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_59 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_60 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_61 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_62 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_63 : OUT STD_LOGIC_VECTOR (15 downto 0) );
    end component;


    component relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0) );
    end component;


    component relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s IS
    port (
        ap_ready : OUT STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_5_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_6_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_7_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_8_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_9_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_10_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_11_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_12_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_13_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_14_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_15_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_16_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_17_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_18_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_19_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_20_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_21_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_22_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_23_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_24_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_25_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_26_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_27_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_28_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_29_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_30_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_31_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_5 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_6 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_7 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_8 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_9 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_10 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_11 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_12 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_13 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_14 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_15 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_16 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_17 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_18 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_19 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_20 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_21 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_22 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_23 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_24 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_25 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_26 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_27 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_28 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_29 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_30 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_31 : OUT STD_LOGIC_VECTOR (15 downto 0) );
    end component;


    component softmax_latency_ap_fixed_ap_fixed_softmax_config13_s IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        ap_start : IN STD_LOGIC;
        ap_done : OUT STD_LOGIC;
        ap_idle : OUT STD_LOGIC;
        ap_ready : OUT STD_LOGIC;
        ap_ce : IN STD_LOGIC;
        data_0_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_1_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_2_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_3_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        data_4_V_read : IN STD_LOGIC_VECTOR (15 downto 0);
        ap_return_0 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_1 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_2 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_3 : OUT STD_LOGIC_VECTOR (15 downto 0);
        ap_return_4 : OUT STD_LOGIC_VECTOR (15 downto 0) );
    end component;



begin
    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_0_V_read => layer4_out_0_V_reg_1821,
        data_1_V_read => layer4_out_1_V_reg_1826,
        data_2_V_read => layer4_out_2_V_reg_1831,
        data_3_V_read => layer4_out_3_V_reg_1836,
        data_4_V_read => layer4_out_4_V_reg_1841,
        data_5_V_read => layer4_out_5_V_reg_1846,
        data_6_V_read => layer4_out_6_V_reg_1851,
        data_7_V_read => layer4_out_7_V_reg_1856,
        data_8_V_read => layer4_out_8_V_reg_1861,
        data_9_V_read => layer4_out_9_V_reg_1866,
        data_10_V_read => layer4_out_10_V_reg_1871,
        data_11_V_read => layer4_out_11_V_reg_1876,
        data_12_V_read => layer4_out_12_V_reg_1881,
        data_13_V_read => layer4_out_13_V_reg_1886,
        data_14_V_read => layer4_out_14_V_reg_1891,
        data_15_V_read => layer4_out_15_V_reg_1896,
        data_16_V_read => layer4_out_16_V_reg_1901,
        data_17_V_read => layer4_out_17_V_reg_1906,
        data_18_V_read => layer4_out_18_V_reg_1911,
        data_19_V_read => layer4_out_19_V_reg_1916,
        data_20_V_read => layer4_out_20_V_reg_1921,
        data_21_V_read => layer4_out_21_V_reg_1926,
        data_22_V_read => layer4_out_22_V_reg_1931,
        data_23_V_read => layer4_out_23_V_reg_1936,
        data_24_V_read => layer4_out_24_V_reg_1941,
        data_25_V_read => layer4_out_25_V_reg_1946,
        data_26_V_read => layer4_out_26_V_reg_1951,
        data_27_V_read => layer4_out_27_V_reg_1956,
        data_28_V_read => layer4_out_28_V_reg_1961,
        data_29_V_read => layer4_out_29_V_reg_1966,
        data_30_V_read => layer4_out_30_V_reg_1971,
        data_31_V_read => layer4_out_31_V_reg_1976,
        data_32_V_read => layer4_out_32_V_reg_1981,
        data_33_V_read => layer4_out_33_V_reg_1986,
        data_34_V_read => layer4_out_34_V_reg_1991,
        data_35_V_read => layer4_out_35_V_reg_1996,
        data_36_V_read => layer4_out_36_V_reg_2001,
        data_37_V_read => layer4_out_37_V_reg_2006,
        data_38_V_read => layer4_out_38_V_reg_2011,
        data_39_V_read => layer4_out_39_V_reg_2016,
        data_40_V_read => layer4_out_40_V_reg_2021,
        data_41_V_read => layer4_out_41_V_reg_2026,
        data_42_V_read => layer4_out_42_V_reg_2031,
        data_43_V_read => layer4_out_43_V_reg_2036,
        data_44_V_read => layer4_out_44_V_reg_2041,
        data_45_V_read => layer4_out_45_V_reg_2046,
        data_46_V_read => layer4_out_46_V_reg_2051,
        data_47_V_read => layer4_out_47_V_reg_2056,
        data_48_V_read => layer4_out_48_V_reg_2061,
        data_49_V_read => layer4_out_49_V_reg_2066,
        data_50_V_read => layer4_out_50_V_reg_2071,
        data_51_V_read => layer4_out_51_V_reg_2076,
        data_52_V_read => layer4_out_52_V_reg_2081,
        data_53_V_read => layer4_out_53_V_reg_2086,
        data_54_V_read => layer4_out_54_V_reg_2091,
        data_55_V_read => layer4_out_55_V_reg_2096,
        data_56_V_read => layer4_out_56_V_reg_2101,
        data_57_V_read => layer4_out_57_V_reg_2106,
        data_58_V_read => layer4_out_58_V_reg_2111,
        data_59_V_read => layer4_out_59_V_reg_2116,
        data_60_V_read => layer4_out_60_V_reg_2121,
        data_61_V_read => layer4_out_61_V_reg_2126,
        data_62_V_read => layer4_out_62_V_reg_2131,
        data_63_V_read => layer4_out_63_V_reg_2136,
        ap_return_0 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_0,
        ap_return_1 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_1,
        ap_return_2 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_2,
        ap_return_3 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_3,
        ap_return_4 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_4,
        ap_return_5 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_5,
        ap_return_6 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_6,
        ap_return_7 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_7,
        ap_return_8 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_8,
        ap_return_9 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_9,
        ap_return_10 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_10,
        ap_return_11 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_11,
        ap_return_12 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_12,
        ap_return_13 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_13,
        ap_return_14 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_14,
        ap_return_15 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_15,
        ap_return_16 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_16,
        ap_return_17 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_17,
        ap_return_18 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_18,
        ap_return_19 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_19,
        ap_return_20 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_20,
        ap_return_21 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_21,
        ap_return_22 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_22,
        ap_return_23 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_23,
        ap_return_24 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_24,
        ap_return_25 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_25,
        ap_return_26 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_26,
        ap_return_27 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_27,
        ap_return_28 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_28,
        ap_return_29 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_29,
        ap_return_30 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_30,
        ap_return_31 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_31,
        ap_ce => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_ce);

    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_V_read => fc1_input_V_in_sig,
        ap_return_0 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_0,
        ap_return_1 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_1,
        ap_return_2 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_2,
        ap_return_3 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_3,
        ap_return_4 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_4,
        ap_return_5 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_5,
        ap_return_6 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_6,
        ap_return_7 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_7,
        ap_return_8 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_8,
        ap_return_9 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_9,
        ap_return_10 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_10,
        ap_return_11 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_11,
        ap_return_12 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_12,
        ap_return_13 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_13,
        ap_return_14 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_14,
        ap_return_15 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_15,
        ap_return_16 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_16,
        ap_return_17 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_17,
        ap_return_18 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_18,
        ap_return_19 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_19,
        ap_return_20 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_20,
        ap_return_21 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_21,
        ap_return_22 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_22,
        ap_return_23 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_23,
        ap_return_24 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_24,
        ap_return_25 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_25,
        ap_return_26 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_26,
        ap_return_27 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_27,
        ap_return_28 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_28,
        ap_return_29 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_29,
        ap_return_30 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_30,
        ap_return_31 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_31,
        ap_return_32 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_32,
        ap_return_33 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_33,
        ap_return_34 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_34,
        ap_return_35 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_35,
        ap_return_36 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_36,
        ap_return_37 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_37,
        ap_return_38 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_38,
        ap_return_39 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_39,
        ap_return_40 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_40,
        ap_return_41 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_41,
        ap_return_42 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_42,
        ap_return_43 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_43,
        ap_return_44 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_44,
        ap_return_45 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_45,
        ap_return_46 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_46,
        ap_return_47 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_47,
        ap_return_48 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_48,
        ap_return_49 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_49,
        ap_return_50 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_50,
        ap_return_51 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_51,
        ap_return_52 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_52,
        ap_return_53 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_53,
        ap_return_54 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_54,
        ap_return_55 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_55,
        ap_return_56 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_56,
        ap_return_57 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_57,
        ap_return_58 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_58,
        ap_return_59 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_59,
        ap_return_60 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_60,
        ap_return_61 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_61,
        ap_return_62 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_62,
        ap_return_63 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_63,
        ap_ce => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_ce);

    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197 : component dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_0_V_read => layer7_out_0_V_reg_2301,
        data_1_V_read => layer7_out_1_V_reg_2306,
        data_2_V_read => layer7_out_2_V_reg_2311,
        data_3_V_read => layer7_out_3_V_reg_2316,
        data_4_V_read => layer7_out_4_V_reg_2321,
        data_5_V_read => layer7_out_5_V_reg_2326,
        data_6_V_read => layer7_out_6_V_reg_2331,
        data_7_V_read => layer7_out_7_V_reg_2336,
        data_8_V_read => layer7_out_8_V_reg_2341,
        data_9_V_read => layer7_out_9_V_reg_2346,
        data_10_V_read => layer7_out_10_V_reg_2351,
        data_11_V_read => layer7_out_11_V_reg_2356,
        data_12_V_read => layer7_out_12_V_reg_2361,
        data_13_V_read => layer7_out_13_V_reg_2366,
        data_14_V_read => layer7_out_14_V_reg_2371,
        data_15_V_read => layer7_out_15_V_reg_2376,
        data_16_V_read => layer7_out_16_V_reg_2381,
        data_17_V_read => layer7_out_17_V_reg_2386,
        data_18_V_read => layer7_out_18_V_reg_2391,
        data_19_V_read => layer7_out_19_V_reg_2396,
        data_20_V_read => layer7_out_20_V_reg_2401,
        data_21_V_read => layer7_out_21_V_reg_2406,
        data_22_V_read => layer7_out_22_V_reg_2411,
        data_23_V_read => layer7_out_23_V_reg_2416,
        data_24_V_read => layer7_out_24_V_reg_2421,
        data_25_V_read => layer7_out_25_V_reg_2426,
        data_26_V_read => layer7_out_26_V_reg_2431,
        data_27_V_read => layer7_out_27_V_reg_2436,
        data_28_V_read => layer7_out_28_V_reg_2441,
        data_29_V_read => layer7_out_29_V_reg_2446,
        data_30_V_read => layer7_out_30_V_reg_2451,
        data_31_V_read => layer7_out_31_V_reg_2456,
        ap_return_0 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_0,
        ap_return_1 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_1,
        ap_return_2 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_2,
        ap_return_3 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_3,
        ap_return_4 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_4,
        ap_return_5 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_5,
        ap_return_6 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_6,
        ap_return_7 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_7,
        ap_return_8 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_8,
        ap_return_9 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_9,
        ap_return_10 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_10,
        ap_return_11 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_11,
        ap_return_12 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_12,
        ap_return_13 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_13,
        ap_return_14 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_14,
        ap_return_15 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_15,
        ap_return_16 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_16,
        ap_return_17 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_17,
        ap_return_18 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_18,
        ap_return_19 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_19,
        ap_return_20 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_20,
        ap_return_21 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_21,
        ap_return_22 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_22,
        ap_return_23 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_23,
        ap_return_24 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_24,
        ap_return_25 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_25,
        ap_return_26 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_26,
        ap_return_27 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_27,
        ap_return_28 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_28,
        ap_return_29 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_29,
        ap_return_30 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_30,
        ap_return_31 => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_31,
        ap_ce => grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_ce);

    grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233 : component dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        data_0_V_read => layer10_out_0_V_reg_2621,
        data_1_V_read => layer10_out_1_V_reg_2626,
        data_2_V_read => layer10_out_2_V_reg_2631,
        data_3_V_read => layer10_out_3_V_reg_2636,
        data_4_V_read => layer10_out_4_V_reg_2641,
        data_5_V_read => layer10_out_5_V_reg_2646,
        data_6_V_read => layer10_out_6_V_reg_2651,
        data_7_V_read => layer10_out_7_V_reg_2656,
        data_8_V_read => layer10_out_8_V_reg_2661,
        data_9_V_read => layer10_out_9_V_reg_2666,
        data_10_V_read => layer10_out_10_V_reg_2671,
        data_11_V_read => layer10_out_11_V_reg_2676,
        data_12_V_read => layer10_out_12_V_reg_2681,
        data_13_V_read => layer10_out_13_V_reg_2686,
        data_14_V_read => layer10_out_14_V_reg_2691,
        data_15_V_read => layer10_out_15_V_reg_2696,
        data_16_V_read => layer10_out_16_V_reg_2701,
        data_17_V_read => layer10_out_17_V_reg_2706,
        data_18_V_read => layer10_out_18_V_reg_2711,
        data_19_V_read => layer10_out_19_V_reg_2716,
        data_20_V_read => layer10_out_20_V_reg_2721,
        data_21_V_read => layer10_out_21_V_reg_2726,
        data_22_V_read => layer10_out_22_V_reg_2731,
        data_23_V_read => layer10_out_23_V_reg_2736,
        data_24_V_read => layer10_out_24_V_reg_2741,
        data_25_V_read => layer10_out_25_V_reg_2746,
        data_26_V_read => layer10_out_26_V_reg_2751,
        data_27_V_read => layer10_out_27_V_reg_2756,
        data_28_V_read => layer10_out_28_V_reg_2761,
        data_29_V_read => layer10_out_29_V_reg_2766,
        data_30_V_read => layer10_out_30_V_reg_2771,
        data_31_V_read => layer10_out_31_V_reg_2776,
        ap_return_0 => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_0,
        ap_return_1 => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_1,
        ap_return_2 => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_2,
        ap_return_3 => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_3,
        ap_return_4 => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_4,
        ap_ce => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_ce);

    call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269 : component relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s
    port map (
        ap_ready => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_ready,
        data_0_V_read => layer2_out_0_V_reg_1501,
        data_1_V_read => layer2_out_1_V_reg_1506,
        data_2_V_read => layer2_out_2_V_reg_1511,
        data_3_V_read => layer2_out_3_V_reg_1516,
        data_4_V_read => layer2_out_4_V_reg_1521,
        data_5_V_read => layer2_out_5_V_reg_1526,
        data_6_V_read => layer2_out_6_V_reg_1531,
        data_7_V_read => layer2_out_7_V_reg_1536,
        data_8_V_read => layer2_out_8_V_reg_1541,
        data_9_V_read => layer2_out_9_V_reg_1546,
        data_10_V_read => layer2_out_10_V_reg_1551,
        data_11_V_read => layer2_out_11_V_reg_1556,
        data_12_V_read => layer2_out_12_V_reg_1561,
        data_13_V_read => layer2_out_13_V_reg_1566,
        data_14_V_read => layer2_out_14_V_reg_1571,
        data_15_V_read => layer2_out_15_V_reg_1576,
        data_16_V_read => layer2_out_16_V_reg_1581,
        data_17_V_read => layer2_out_17_V_reg_1586,
        data_18_V_read => layer2_out_18_V_reg_1591,
        data_19_V_read => layer2_out_19_V_reg_1596,
        data_20_V_read => layer2_out_20_V_reg_1601,
        data_21_V_read => layer2_out_21_V_reg_1606,
        data_22_V_read => layer2_out_22_V_reg_1611,
        data_23_V_read => layer2_out_23_V_reg_1616,
        data_24_V_read => layer2_out_24_V_reg_1621,
        data_25_V_read => layer2_out_25_V_reg_1626,
        data_26_V_read => layer2_out_26_V_reg_1631,
        data_27_V_read => layer2_out_27_V_reg_1636,
        data_28_V_read => layer2_out_28_V_reg_1641,
        data_29_V_read => layer2_out_29_V_reg_1646,
        data_30_V_read => layer2_out_30_V_reg_1651,
        data_31_V_read => layer2_out_31_V_reg_1656,
        data_32_V_read => layer2_out_32_V_reg_1661,
        data_33_V_read => layer2_out_33_V_reg_1666,
        data_34_V_read => layer2_out_34_V_reg_1671,
        data_35_V_read => layer2_out_35_V_reg_1676,
        data_36_V_read => layer2_out_36_V_reg_1681,
        data_37_V_read => layer2_out_37_V_reg_1686,
        data_38_V_read => layer2_out_38_V_reg_1691,
        data_39_V_read => layer2_out_39_V_reg_1696,
        data_40_V_read => layer2_out_40_V_reg_1701,
        data_41_V_read => layer2_out_41_V_reg_1706,
        data_42_V_read => layer2_out_42_V_reg_1711,
        data_43_V_read => layer2_out_43_V_reg_1716,
        data_44_V_read => layer2_out_44_V_reg_1721,
        data_45_V_read => layer2_out_45_V_reg_1726,
        data_46_V_read => layer2_out_46_V_reg_1731,
        data_47_V_read => layer2_out_47_V_reg_1736,
        data_48_V_read => layer2_out_48_V_reg_1741,
        data_49_V_read => layer2_out_49_V_reg_1746,
        data_50_V_read => layer2_out_50_V_reg_1751,
        data_51_V_read => layer2_out_51_V_reg_1756,
        data_52_V_read => layer2_out_52_V_reg_1761,
        data_53_V_read => layer2_out_53_V_reg_1766,
        data_54_V_read => layer2_out_54_V_reg_1771,
        data_55_V_read => layer2_out_55_V_reg_1776,
        data_56_V_read => layer2_out_56_V_reg_1781,
        data_57_V_read => layer2_out_57_V_reg_1786,
        data_58_V_read => layer2_out_58_V_reg_1791,
        data_59_V_read => layer2_out_59_V_reg_1796,
        data_60_V_read => layer2_out_60_V_reg_1801,
        data_61_V_read => layer2_out_61_V_reg_1806,
        data_62_V_read => layer2_out_62_V_reg_1811,
        data_63_V_read => layer2_out_63_V_reg_1816,
        ap_return_0 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_0,
        ap_return_1 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_1,
        ap_return_2 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_2,
        ap_return_3 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_3,
        ap_return_4 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_4,
        ap_return_5 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_5,
        ap_return_6 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_6,
        ap_return_7 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_7,
        ap_return_8 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_8,
        ap_return_9 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_9,
        ap_return_10 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_10,
        ap_return_11 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_11,
        ap_return_12 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_12,
        ap_return_13 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_13,
        ap_return_14 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_14,
        ap_return_15 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_15,
        ap_return_16 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_16,
        ap_return_17 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_17,
        ap_return_18 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_18,
        ap_return_19 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_19,
        ap_return_20 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_20,
        ap_return_21 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_21,
        ap_return_22 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_22,
        ap_return_23 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_23,
        ap_return_24 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_24,
        ap_return_25 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_25,
        ap_return_26 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_26,
        ap_return_27 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_27,
        ap_return_28 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_28,
        ap_return_29 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_29,
        ap_return_30 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_30,
        ap_return_31 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_31,
        ap_return_32 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_32,
        ap_return_33 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_33,
        ap_return_34 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_34,
        ap_return_35 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_35,
        ap_return_36 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_36,
        ap_return_37 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_37,
        ap_return_38 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_38,
        ap_return_39 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_39,
        ap_return_40 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_40,
        ap_return_41 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_41,
        ap_return_42 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_42,
        ap_return_43 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_43,
        ap_return_44 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_44,
        ap_return_45 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_45,
        ap_return_46 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_46,
        ap_return_47 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_47,
        ap_return_48 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_48,
        ap_return_49 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_49,
        ap_return_50 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_50,
        ap_return_51 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_51,
        ap_return_52 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_52,
        ap_return_53 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_53,
        ap_return_54 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_54,
        ap_return_55 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_55,
        ap_return_56 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_56,
        ap_return_57 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_57,
        ap_return_58 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_58,
        ap_return_59 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_59,
        ap_return_60 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_60,
        ap_return_61 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_61,
        ap_return_62 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_62,
        ap_return_63 => call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_63);

    call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337 : component relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s
    port map (
        ap_ready => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_ready,
        data_0_V_read => layer5_out_0_V_reg_2141,
        data_1_V_read => layer5_out_1_V_reg_2146,
        data_2_V_read => layer5_out_2_V_reg_2151,
        data_3_V_read => layer5_out_3_V_reg_2156,
        data_4_V_read => layer5_out_4_V_reg_2161,
        data_5_V_read => layer5_out_5_V_reg_2166,
        data_6_V_read => layer5_out_6_V_reg_2171,
        data_7_V_read => layer5_out_7_V_reg_2176,
        data_8_V_read => layer5_out_8_V_reg_2181,
        data_9_V_read => layer5_out_9_V_reg_2186,
        data_10_V_read => layer5_out_10_V_reg_2191,
        data_11_V_read => layer5_out_11_V_reg_2196,
        data_12_V_read => layer5_out_12_V_reg_2201,
        data_13_V_read => layer5_out_13_V_reg_2206,
        data_14_V_read => layer5_out_14_V_reg_2211,
        data_15_V_read => layer5_out_15_V_reg_2216,
        data_16_V_read => layer5_out_16_V_reg_2221,
        data_17_V_read => layer5_out_17_V_reg_2226,
        data_18_V_read => layer5_out_18_V_reg_2231,
        data_19_V_read => layer5_out_19_V_reg_2236,
        data_20_V_read => layer5_out_20_V_reg_2241,
        data_21_V_read => layer5_out_21_V_reg_2246,
        data_22_V_read => layer5_out_22_V_reg_2251,
        data_23_V_read => layer5_out_23_V_reg_2256,
        data_24_V_read => layer5_out_24_V_reg_2261,
        data_25_V_read => layer5_out_25_V_reg_2266,
        data_26_V_read => layer5_out_26_V_reg_2271,
        data_27_V_read => layer5_out_27_V_reg_2276,
        data_28_V_read => layer5_out_28_V_reg_2281,
        data_29_V_read => layer5_out_29_V_reg_2286,
        data_30_V_read => layer5_out_30_V_reg_2291,
        data_31_V_read => layer5_out_31_V_reg_2296,
        ap_return_0 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_0,
        ap_return_1 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_1,
        ap_return_2 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_2,
        ap_return_3 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_3,
        ap_return_4 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_4,
        ap_return_5 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_5,
        ap_return_6 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_6,
        ap_return_7 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_7,
        ap_return_8 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_8,
        ap_return_9 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_9,
        ap_return_10 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_10,
        ap_return_11 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_11,
        ap_return_12 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_12,
        ap_return_13 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_13,
        ap_return_14 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_14,
        ap_return_15 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_15,
        ap_return_16 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_16,
        ap_return_17 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_17,
        ap_return_18 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_18,
        ap_return_19 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_19,
        ap_return_20 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_20,
        ap_return_21 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_21,
        ap_return_22 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_22,
        ap_return_23 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_23,
        ap_return_24 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_24,
        ap_return_25 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_25,
        ap_return_26 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_26,
        ap_return_27 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_27,
        ap_return_28 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_28,
        ap_return_29 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_29,
        ap_return_30 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_30,
        ap_return_31 => call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_31);

    call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373 : component relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s
    port map (
        ap_ready => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_ready,
        data_0_V_read => layer8_out_0_V_reg_2461,
        data_1_V_read => layer8_out_1_V_reg_2466,
        data_2_V_read => layer8_out_2_V_reg_2471,
        data_3_V_read => layer8_out_3_V_reg_2476,
        data_4_V_read => layer8_out_4_V_reg_2481,
        data_5_V_read => layer8_out_5_V_reg_2486,
        data_6_V_read => layer8_out_6_V_reg_2491,
        data_7_V_read => layer8_out_7_V_reg_2496,
        data_8_V_read => layer8_out_8_V_reg_2501,
        data_9_V_read => layer8_out_9_V_reg_2506,
        data_10_V_read => layer8_out_10_V_reg_2511,
        data_11_V_read => layer8_out_11_V_reg_2516,
        data_12_V_read => layer8_out_12_V_reg_2521,
        data_13_V_read => layer8_out_13_V_reg_2526,
        data_14_V_read => layer8_out_14_V_reg_2531,
        data_15_V_read => layer8_out_15_V_reg_2536,
        data_16_V_read => layer8_out_16_V_reg_2541,
        data_17_V_read => layer8_out_17_V_reg_2546,
        data_18_V_read => layer8_out_18_V_reg_2551,
        data_19_V_read => layer8_out_19_V_reg_2556,
        data_20_V_read => layer8_out_20_V_reg_2561,
        data_21_V_read => layer8_out_21_V_reg_2566,
        data_22_V_read => layer8_out_22_V_reg_2571,
        data_23_V_read => layer8_out_23_V_reg_2576,
        data_24_V_read => layer8_out_24_V_reg_2581,
        data_25_V_read => layer8_out_25_V_reg_2586,
        data_26_V_read => layer8_out_26_V_reg_2591,
        data_27_V_read => layer8_out_27_V_reg_2596,
        data_28_V_read => layer8_out_28_V_reg_2601,
        data_29_V_read => layer8_out_29_V_reg_2606,
        data_30_V_read => layer8_out_30_V_reg_2611,
        data_31_V_read => layer8_out_31_V_reg_2616,
        ap_return_0 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_0,
        ap_return_1 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_1,
        ap_return_2 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_2,
        ap_return_3 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_3,
        ap_return_4 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_4,
        ap_return_5 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_5,
        ap_return_6 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_6,
        ap_return_7 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_7,
        ap_return_8 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_8,
        ap_return_9 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_9,
        ap_return_10 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_10,
        ap_return_11 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_11,
        ap_return_12 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_12,
        ap_return_13 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_13,
        ap_return_14 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_14,
        ap_return_15 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_15,
        ap_return_16 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_16,
        ap_return_17 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_17,
        ap_return_18 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_18,
        ap_return_19 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_19,
        ap_return_20 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_20,
        ap_return_21 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_21,
        ap_return_22 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_22,
        ap_return_23 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_23,
        ap_return_24 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_24,
        ap_return_25 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_25,
        ap_return_26 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_26,
        ap_return_27 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_27,
        ap_return_28 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_28,
        ap_return_29 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_29,
        ap_return_30 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_30,
        ap_return_31 => call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_31);

    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409 : component softmax_latency_ap_fixed_ap_fixed_softmax_config13_s
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        ap_start => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start,
        ap_done => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_done,
        ap_idle => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_idle,
        ap_ready => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_ready,
        ap_ce => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_ce,
        data_0_V_read => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_0,
        data_1_V_read => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_1,
        data_2_V_read => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_2,
        data_3_V_read => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_3,
        data_4_V_read => grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_return_4,
        ap_return_0 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_0,
        ap_return_1 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_1,
        ap_return_2 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_2,
        ap_return_3 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_3,
        ap_return_4 => grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_4);





    ap_CS_fsm_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
            else
                ap_CS_fsm <= ap_NS_fsm;
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter1_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter1 <= ap_const_logic_0;
            else
                if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_subdone))) then 
                    ap_enable_reg_pp0_iter1 <= ap_start;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter10_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter10 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter11_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter11 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter12_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter12 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter13_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter13 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter14_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter14 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter15_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter15 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter16_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter16 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter17_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter17 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter18_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter18 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter19_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter19 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter2_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter2 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter20_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter20 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter21_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter21 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter22_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter22 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter23_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter23 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter24_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter24 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter25_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter25 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter26_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter26 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter27_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter27 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter27 <= ap_enable_reg_pp0_iter26;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter28_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter28 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter28 <= ap_enable_reg_pp0_iter27;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter29_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter29 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter29 <= ap_enable_reg_pp0_iter28;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter3_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter3 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter30_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter30 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter30 <= ap_enable_reg_pp0_iter29;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter31_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter31 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter31 <= ap_enable_reg_pp0_iter30;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter32_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter32 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter32 <= ap_enable_reg_pp0_iter31;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter33_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter33 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter33 <= ap_enable_reg_pp0_iter32;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter34_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter34 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter34 <= ap_enable_reg_pp0_iter33;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter35_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter35 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter35 <= ap_enable_reg_pp0_iter34;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter36_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter36 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter36 <= ap_enable_reg_pp0_iter35;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter37_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter37 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter37 <= ap_enable_reg_pp0_iter36;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter38_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter38 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter38 <= ap_enable_reg_pp0_iter37;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter4_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter4 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter5_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter5 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter6_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter6 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter7_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter7 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter8_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter8 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter9_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_enable_reg_pp0_iter9 <= ap_const_logic_0;
            else
                if ((ap_const_boolean_0 = ap_block_pp0_stage0_subdone)) then 
                    ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
                end if; 
            end if;
        end if;
    end process;


    fc1_input_V_ap_vld_preg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                fc1_input_V_ap_vld_preg <= ap_const_logic_0;
            else
                if (((ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
                    fc1_input_V_ap_vld_preg <= ap_const_logic_0;
                elsif ((not(((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) and (fc1_input_V_ap_vld = ap_const_logic_1))) then 
                    fc1_input_V_ap_vld_preg <= fc1_input_V_ap_vld;
                end if; 
            end if;
        end if;
    end process;


    fc1_input_V_preg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                fc1_input_V_preg <= ap_const_lv256_lc_1;
            else
                if ((not(((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) and (fc1_input_V_ap_vld = ap_const_logic_1))) then 
                    fc1_input_V_preg <= fc1_input_V;
                end if; 
            end if;
        end if;
    end process;


    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start_reg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start_reg <= ap_const_logic_0;
            else
                if (((ap_enable_reg_pp0_iter30 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
                    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start_reg <= ap_const_logic_1;
                elsif ((grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_ready = ap_const_logic_1)) then 
                    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start_reg <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;

    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_const_boolean_0 = ap_block_pp0_stage0_11001)) then
                layer10_out_0_V_reg_2621 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_0;
                layer10_out_10_V_reg_2671 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_10;
                layer10_out_11_V_reg_2676 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_11;
                layer10_out_12_V_reg_2681 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_12;
                layer10_out_13_V_reg_2686 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_13;
                layer10_out_14_V_reg_2691 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_14;
                layer10_out_15_V_reg_2696 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_15;
                layer10_out_16_V_reg_2701 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_16;
                layer10_out_17_V_reg_2706 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_17;
                layer10_out_18_V_reg_2711 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_18;
                layer10_out_19_V_reg_2716 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_19;
                layer10_out_1_V_reg_2626 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_1;
                layer10_out_20_V_reg_2721 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_20;
                layer10_out_21_V_reg_2726 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_21;
                layer10_out_22_V_reg_2731 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_22;
                layer10_out_23_V_reg_2736 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_23;
                layer10_out_24_V_reg_2741 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_24;
                layer10_out_25_V_reg_2746 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_25;
                layer10_out_26_V_reg_2751 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_26;
                layer10_out_27_V_reg_2756 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_27;
                layer10_out_28_V_reg_2761 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_28;
                layer10_out_29_V_reg_2766 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_29;
                layer10_out_2_V_reg_2631 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_2;
                layer10_out_30_V_reg_2771 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_30;
                layer10_out_31_V_reg_2776 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_31;
                layer10_out_3_V_reg_2636 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_3;
                layer10_out_4_V_reg_2641 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_4;
                layer10_out_5_V_reg_2646 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_5;
                layer10_out_6_V_reg_2651 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_6;
                layer10_out_7_V_reg_2656 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_7;
                layer10_out_8_V_reg_2661 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_8;
                layer10_out_9_V_reg_2666 <= call_ret5_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config10_s_fu_373_ap_return_9;
                layer2_out_0_V_reg_1501 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_0;
                layer2_out_10_V_reg_1551 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_10;
                layer2_out_11_V_reg_1556 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_11;
                layer2_out_12_V_reg_1561 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_12;
                layer2_out_13_V_reg_1566 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_13;
                layer2_out_14_V_reg_1571 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_14;
                layer2_out_15_V_reg_1576 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_15;
                layer2_out_16_V_reg_1581 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_16;
                layer2_out_17_V_reg_1586 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_17;
                layer2_out_18_V_reg_1591 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_18;
                layer2_out_19_V_reg_1596 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_19;
                layer2_out_1_V_reg_1506 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_1;
                layer2_out_20_V_reg_1601 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_20;
                layer2_out_21_V_reg_1606 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_21;
                layer2_out_22_V_reg_1611 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_22;
                layer2_out_23_V_reg_1616 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_23;
                layer2_out_24_V_reg_1621 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_24;
                layer2_out_25_V_reg_1626 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_25;
                layer2_out_26_V_reg_1631 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_26;
                layer2_out_27_V_reg_1636 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_27;
                layer2_out_28_V_reg_1641 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_28;
                layer2_out_29_V_reg_1646 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_29;
                layer2_out_2_V_reg_1511 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_2;
                layer2_out_30_V_reg_1651 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_30;
                layer2_out_31_V_reg_1656 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_31;
                layer2_out_32_V_reg_1661 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_32;
                layer2_out_33_V_reg_1666 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_33;
                layer2_out_34_V_reg_1671 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_34;
                layer2_out_35_V_reg_1676 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_35;
                layer2_out_36_V_reg_1681 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_36;
                layer2_out_37_V_reg_1686 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_37;
                layer2_out_38_V_reg_1691 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_38;
                layer2_out_39_V_reg_1696 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_39;
                layer2_out_3_V_reg_1516 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_3;
                layer2_out_40_V_reg_1701 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_40;
                layer2_out_41_V_reg_1706 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_41;
                layer2_out_42_V_reg_1711 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_42;
                layer2_out_43_V_reg_1716 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_43;
                layer2_out_44_V_reg_1721 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_44;
                layer2_out_45_V_reg_1726 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_45;
                layer2_out_46_V_reg_1731 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_46;
                layer2_out_47_V_reg_1736 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_47;
                layer2_out_48_V_reg_1741 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_48;
                layer2_out_49_V_reg_1746 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_49;
                layer2_out_4_V_reg_1521 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_4;
                layer2_out_50_V_reg_1751 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_50;
                layer2_out_51_V_reg_1756 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_51;
                layer2_out_52_V_reg_1761 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_52;
                layer2_out_53_V_reg_1766 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_53;
                layer2_out_54_V_reg_1771 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_54;
                layer2_out_55_V_reg_1776 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_55;
                layer2_out_56_V_reg_1781 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_56;
                layer2_out_57_V_reg_1786 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_57;
                layer2_out_58_V_reg_1791 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_58;
                layer2_out_59_V_reg_1796 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_59;
                layer2_out_5_V_reg_1526 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_5;
                layer2_out_60_V_reg_1801 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_60;
                layer2_out_61_V_reg_1806 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_61;
                layer2_out_62_V_reg_1811 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_62;
                layer2_out_63_V_reg_1816 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_63;
                layer2_out_6_V_reg_1531 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_6;
                layer2_out_7_V_reg_1536 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_7;
                layer2_out_8_V_reg_1541 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_8;
                layer2_out_9_V_reg_1546 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_return_9;
                layer4_out_0_V_reg_1821 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_0;
                layer4_out_10_V_reg_1871 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_10;
                layer4_out_11_V_reg_1876 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_11;
                layer4_out_12_V_reg_1881 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_12;
                layer4_out_13_V_reg_1886 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_13;
                layer4_out_14_V_reg_1891 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_14;
                layer4_out_15_V_reg_1896 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_15;
                layer4_out_16_V_reg_1901 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_16;
                layer4_out_17_V_reg_1906 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_17;
                layer4_out_18_V_reg_1911 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_18;
                layer4_out_19_V_reg_1916 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_19;
                layer4_out_1_V_reg_1826 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_1;
                layer4_out_20_V_reg_1921 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_20;
                layer4_out_21_V_reg_1926 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_21;
                layer4_out_22_V_reg_1931 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_22;
                layer4_out_23_V_reg_1936 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_23;
                layer4_out_24_V_reg_1941 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_24;
                layer4_out_25_V_reg_1946 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_25;
                layer4_out_26_V_reg_1951 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_26;
                layer4_out_27_V_reg_1956 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_27;
                layer4_out_28_V_reg_1961 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_28;
                layer4_out_29_V_reg_1966 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_29;
                layer4_out_2_V_reg_1831 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_2;
                layer4_out_30_V_reg_1971 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_30;
                layer4_out_31_V_reg_1976 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_31;
                layer4_out_32_V_reg_1981 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_32;
                layer4_out_33_V_reg_1986 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_33;
                layer4_out_34_V_reg_1991 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_34;
                layer4_out_35_V_reg_1996 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_35;
                layer4_out_36_V_reg_2001 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_36;
                layer4_out_37_V_reg_2006 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_37;
                layer4_out_38_V_reg_2011 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_38;
                layer4_out_39_V_reg_2016 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_39;
                layer4_out_3_V_reg_1836 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_3;
                layer4_out_40_V_reg_2021 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_40;
                layer4_out_41_V_reg_2026 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_41;
                layer4_out_42_V_reg_2031 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_42;
                layer4_out_43_V_reg_2036 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_43;
                layer4_out_44_V_reg_2041 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_44;
                layer4_out_45_V_reg_2046 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_45;
                layer4_out_46_V_reg_2051 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_46;
                layer4_out_47_V_reg_2056 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_47;
                layer4_out_48_V_reg_2061 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_48;
                layer4_out_49_V_reg_2066 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_49;
                layer4_out_4_V_reg_1841 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_4;
                layer4_out_50_V_reg_2071 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_50;
                layer4_out_51_V_reg_2076 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_51;
                layer4_out_52_V_reg_2081 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_52;
                layer4_out_53_V_reg_2086 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_53;
                layer4_out_54_V_reg_2091 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_54;
                layer4_out_55_V_reg_2096 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_55;
                layer4_out_56_V_reg_2101 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_56;
                layer4_out_57_V_reg_2106 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_57;
                layer4_out_58_V_reg_2111 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_58;
                layer4_out_59_V_reg_2116 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_59;
                layer4_out_5_V_reg_1846 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_5;
                layer4_out_60_V_reg_2121 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_60;
                layer4_out_61_V_reg_2126 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_61;
                layer4_out_62_V_reg_2131 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_62;
                layer4_out_63_V_reg_2136 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_63;
                layer4_out_6_V_reg_1851 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_6;
                layer4_out_7_V_reg_1856 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_7;
                layer4_out_8_V_reg_1861 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_8;
                layer4_out_9_V_reg_1866 <= call_ret1_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config4_s_fu_269_ap_return_9;
                layer5_out_0_V_reg_2141 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_0;
                layer5_out_10_V_reg_2191 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_10;
                layer5_out_11_V_reg_2196 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_11;
                layer5_out_12_V_reg_2201 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_12;
                layer5_out_13_V_reg_2206 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_13;
                layer5_out_14_V_reg_2211 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_14;
                layer5_out_15_V_reg_2216 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_15;
                layer5_out_16_V_reg_2221 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_16;
                layer5_out_17_V_reg_2226 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_17;
                layer5_out_18_V_reg_2231 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_18;
                layer5_out_19_V_reg_2236 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_19;
                layer5_out_1_V_reg_2146 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_1;
                layer5_out_20_V_reg_2241 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_20;
                layer5_out_21_V_reg_2246 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_21;
                layer5_out_22_V_reg_2251 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_22;
                layer5_out_23_V_reg_2256 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_23;
                layer5_out_24_V_reg_2261 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_24;
                layer5_out_25_V_reg_2266 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_25;
                layer5_out_26_V_reg_2271 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_26;
                layer5_out_27_V_reg_2276 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_27;
                layer5_out_28_V_reg_2281 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_28;
                layer5_out_29_V_reg_2286 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_29;
                layer5_out_2_V_reg_2151 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_2;
                layer5_out_30_V_reg_2291 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_30;
                layer5_out_31_V_reg_2296 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_31;
                layer5_out_3_V_reg_2156 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_3;
                layer5_out_4_V_reg_2161 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_4;
                layer5_out_5_V_reg_2166 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_5;
                layer5_out_6_V_reg_2171 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_6;
                layer5_out_7_V_reg_2176 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_7;
                layer5_out_8_V_reg_2181 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_8;
                layer5_out_9_V_reg_2186 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_return_9;
                layer7_out_0_V_reg_2301 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_0;
                layer7_out_10_V_reg_2351 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_10;
                layer7_out_11_V_reg_2356 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_11;
                layer7_out_12_V_reg_2361 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_12;
                layer7_out_13_V_reg_2366 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_13;
                layer7_out_14_V_reg_2371 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_14;
                layer7_out_15_V_reg_2376 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_15;
                layer7_out_16_V_reg_2381 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_16;
                layer7_out_17_V_reg_2386 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_17;
                layer7_out_18_V_reg_2391 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_18;
                layer7_out_19_V_reg_2396 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_19;
                layer7_out_1_V_reg_2306 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_1;
                layer7_out_20_V_reg_2401 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_20;
                layer7_out_21_V_reg_2406 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_21;
                layer7_out_22_V_reg_2411 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_22;
                layer7_out_23_V_reg_2416 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_23;
                layer7_out_24_V_reg_2421 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_24;
                layer7_out_25_V_reg_2426 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_25;
                layer7_out_26_V_reg_2431 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_26;
                layer7_out_27_V_reg_2436 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_27;
                layer7_out_28_V_reg_2441 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_28;
                layer7_out_29_V_reg_2446 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_29;
                layer7_out_2_V_reg_2311 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_2;
                layer7_out_30_V_reg_2451 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_30;
                layer7_out_31_V_reg_2456 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_31;
                layer7_out_3_V_reg_2316 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_3;
                layer7_out_4_V_reg_2321 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_4;
                layer7_out_5_V_reg_2326 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_5;
                layer7_out_6_V_reg_2331 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_6;
                layer7_out_7_V_reg_2336 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_7;
                layer7_out_8_V_reg_2341 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_8;
                layer7_out_9_V_reg_2346 <= call_ret3_relu_ap_fixed_ap_fixed_16_6_5_3_0_relu_config7_s_fu_337_ap_return_9;
                layer8_out_0_V_reg_2461 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_0;
                layer8_out_10_V_reg_2511 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_10;
                layer8_out_11_V_reg_2516 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_11;
                layer8_out_12_V_reg_2521 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_12;
                layer8_out_13_V_reg_2526 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_13;
                layer8_out_14_V_reg_2531 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_14;
                layer8_out_15_V_reg_2536 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_15;
                layer8_out_16_V_reg_2541 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_16;
                layer8_out_17_V_reg_2546 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_17;
                layer8_out_18_V_reg_2551 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_18;
                layer8_out_19_V_reg_2556 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_19;
                layer8_out_1_V_reg_2466 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_1;
                layer8_out_20_V_reg_2561 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_20;
                layer8_out_21_V_reg_2566 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_21;
                layer8_out_22_V_reg_2571 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_22;
                layer8_out_23_V_reg_2576 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_23;
                layer8_out_24_V_reg_2581 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_24;
                layer8_out_25_V_reg_2586 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_25;
                layer8_out_26_V_reg_2591 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_26;
                layer8_out_27_V_reg_2596 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_27;
                layer8_out_28_V_reg_2601 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_28;
                layer8_out_29_V_reg_2606 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_29;
                layer8_out_2_V_reg_2471 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_2;
                layer8_out_30_V_reg_2611 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_30;
                layer8_out_31_V_reg_2616 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_31;
                layer8_out_3_V_reg_2476 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_3;
                layer8_out_4_V_reg_2481 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_4;
                layer8_out_5_V_reg_2486 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_5;
                layer8_out_6_V_reg_2491 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_6;
                layer8_out_7_V_reg_2496 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_7;
                layer8_out_8_V_reg_2501 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_8;
                layer8_out_9_V_reg_2506 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_return_9;
            end if;
        end if;
    end process;

    ap_NS_fsm_assign_proc : process (ap_CS_fsm, ap_block_pp0_stage0_subdone, ap_reset_idle_pp0)
    begin
        case ap_CS_fsm is
            when ap_ST_fsm_pp0_stage0 => 
                ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
            when others =>  
                ap_NS_fsm <= "X";
        end case;
    end process;
    ap_CS_fsm_pp0_stage0 <= ap_CS_fsm(0);
        ap_block_pp0_stage0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage0_01001_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_01001 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp177_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp177 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp250_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp250 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp322_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp322 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp334_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp334 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_11001_ignoreCallOp41_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_11001_ignoreCallOp41 <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;


    ap_block_pp0_stage0_subdone_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_pp0_stage0_subdone <= ((ap_start = ap_const_logic_1) and ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0)));
    end process;

        ap_block_state10_pp0_stage0_iter9 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state10_pp0_stage0_iter9_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state10_pp0_stage0_iter9_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state10_pp0_stage0_iter9_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state10_pp0_stage0_iter9_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state10_pp0_stage0_iter9_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state11_pp0_stage0_iter10_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state12_pp0_stage0_iter11 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state12_pp0_stage0_iter11_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state12_pp0_stage0_iter11_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state12_pp0_stage0_iter11_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state12_pp0_stage0_iter11_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state12_pp0_stage0_iter11_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state13_pp0_stage0_iter12 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state13_pp0_stage0_iter12_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state13_pp0_stage0_iter12_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state13_pp0_stage0_iter12_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state13_pp0_stage0_iter12_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state13_pp0_stage0_iter12_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state14_pp0_stage0_iter13 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state14_pp0_stage0_iter13_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state14_pp0_stage0_iter13_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state14_pp0_stage0_iter13_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state14_pp0_stage0_iter13_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state14_pp0_stage0_iter13_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state15_pp0_stage0_iter14 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state15_pp0_stage0_iter14_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state15_pp0_stage0_iter14_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state15_pp0_stage0_iter14_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state15_pp0_stage0_iter14_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state15_pp0_stage0_iter14_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state16_pp0_stage0_iter15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state16_pp0_stage0_iter15_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state16_pp0_stage0_iter15_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state16_pp0_stage0_iter15_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state16_pp0_stage0_iter15_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state16_pp0_stage0_iter15_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state17_pp0_stage0_iter16 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state17_pp0_stage0_iter16_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state17_pp0_stage0_iter16_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state17_pp0_stage0_iter16_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state17_pp0_stage0_iter16_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state17_pp0_stage0_iter16_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state18_pp0_stage0_iter17 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state18_pp0_stage0_iter17_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state18_pp0_stage0_iter17_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state18_pp0_stage0_iter17_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state18_pp0_stage0_iter17_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state18_pp0_stage0_iter17_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state19_pp0_stage0_iter18 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state19_pp0_stage0_iter18_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state19_pp0_stage0_iter18_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state19_pp0_stage0_iter18_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state19_pp0_stage0_iter18_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state19_pp0_stage0_iter18_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state1_pp0_stage0_iter0_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call145_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call145 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call15_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call15 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call211_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call211 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call277_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call277 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;


    ap_block_state1_pp0_stage0_iter0_ignore_call283_assign_proc : process(ap_start, fc1_input_V_ap_vld_in_sig)
    begin
                ap_block_state1_pp0_stage0_iter0_ignore_call283 <= ((ap_start = ap_const_logic_0) or (fc1_input_V_ap_vld_in_sig = ap_const_logic_0));
    end process;

        ap_block_state20_pp0_stage0_iter19 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state20_pp0_stage0_iter19_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state20_pp0_stage0_iter19_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state20_pp0_stage0_iter19_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state20_pp0_stage0_iter19_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state20_pp0_stage0_iter19_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state21_pp0_stage0_iter20 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state21_pp0_stage0_iter20_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state21_pp0_stage0_iter20_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state21_pp0_stage0_iter20_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state21_pp0_stage0_iter20_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state21_pp0_stage0_iter20_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state22_pp0_stage0_iter21 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state22_pp0_stage0_iter21_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state22_pp0_stage0_iter21_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state22_pp0_stage0_iter21_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state22_pp0_stage0_iter21_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state22_pp0_stage0_iter21_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state23_pp0_stage0_iter22 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state23_pp0_stage0_iter22_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state23_pp0_stage0_iter22_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state23_pp0_stage0_iter22_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state23_pp0_stage0_iter22_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state23_pp0_stage0_iter22_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state24_pp0_stage0_iter23 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state24_pp0_stage0_iter23_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state24_pp0_stage0_iter23_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state24_pp0_stage0_iter23_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state24_pp0_stage0_iter23_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state24_pp0_stage0_iter23_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state25_pp0_stage0_iter24 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state25_pp0_stage0_iter24_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state25_pp0_stage0_iter24_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state25_pp0_stage0_iter24_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state25_pp0_stage0_iter24_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state25_pp0_stage0_iter24_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state26_pp0_stage0_iter25 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state26_pp0_stage0_iter25_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state26_pp0_stage0_iter25_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state26_pp0_stage0_iter25_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state26_pp0_stage0_iter25_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state26_pp0_stage0_iter25_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state27_pp0_stage0_iter26 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state27_pp0_stage0_iter26_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state27_pp0_stage0_iter26_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state27_pp0_stage0_iter26_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state27_pp0_stage0_iter26_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state27_pp0_stage0_iter26_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state28_pp0_stage0_iter27 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state28_pp0_stage0_iter27_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state28_pp0_stage0_iter27_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state28_pp0_stage0_iter27_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state28_pp0_stage0_iter27_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state28_pp0_stage0_iter27_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state29_pp0_stage0_iter28 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state29_pp0_stage0_iter28_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state29_pp0_stage0_iter28_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state29_pp0_stage0_iter28_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state29_pp0_stage0_iter28_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state29_pp0_stage0_iter28_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter1_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state30_pp0_stage0_iter29 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state30_pp0_stage0_iter29_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state30_pp0_stage0_iter29_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state30_pp0_stage0_iter29_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state30_pp0_stage0_iter29_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state30_pp0_stage0_iter29_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state31_pp0_stage0_iter30 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state31_pp0_stage0_iter30_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state31_pp0_stage0_iter30_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state31_pp0_stage0_iter30_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state31_pp0_stage0_iter30_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state31_pp0_stage0_iter30_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state32_pp0_stage0_iter31 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state32_pp0_stage0_iter31_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state32_pp0_stage0_iter31_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state32_pp0_stage0_iter31_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state32_pp0_stage0_iter31_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state32_pp0_stage0_iter31_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state33_pp0_stage0_iter32 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state33_pp0_stage0_iter32_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state33_pp0_stage0_iter32_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state33_pp0_stage0_iter32_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state33_pp0_stage0_iter32_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state33_pp0_stage0_iter32_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state34_pp0_stage0_iter33 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state34_pp0_stage0_iter33_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state34_pp0_stage0_iter33_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state34_pp0_stage0_iter33_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state34_pp0_stage0_iter33_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state34_pp0_stage0_iter33_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state35_pp0_stage0_iter34 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state35_pp0_stage0_iter34_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state35_pp0_stage0_iter34_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state35_pp0_stage0_iter34_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state35_pp0_stage0_iter34_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state35_pp0_stage0_iter34_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state36_pp0_stage0_iter35 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state36_pp0_stage0_iter35_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state36_pp0_stage0_iter35_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state36_pp0_stage0_iter35_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state36_pp0_stage0_iter35_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state36_pp0_stage0_iter35_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state37_pp0_stage0_iter36 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state37_pp0_stage0_iter36_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state37_pp0_stage0_iter36_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state37_pp0_stage0_iter36_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state37_pp0_stage0_iter36_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state37_pp0_stage0_iter36_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state38_pp0_stage0_iter37 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state38_pp0_stage0_iter37_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state38_pp0_stage0_iter37_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state38_pp0_stage0_iter37_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state38_pp0_stage0_iter37_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state38_pp0_stage0_iter37_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state39_pp0_stage0_iter38 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state39_pp0_stage0_iter38_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state39_pp0_stage0_iter38_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state39_pp0_stage0_iter38_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state39_pp0_stage0_iter38_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state39_pp0_stage0_iter38_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state3_pp0_stage0_iter2_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state4_pp0_stage0_iter3_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state5_pp0_stage0_iter4_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage0_iter5_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage0_iter6_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage0_iter7_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call145 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call15 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call211 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call277 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state9_pp0_stage0_iter8_ignore_call283 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_done_assign_proc : process(ap_enable_reg_pp0_iter38, ap_block_pp0_stage0_11001)
    begin
        if (((ap_enable_reg_pp0_iter38 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            ap_done <= ap_const_logic_1;
        else 
            ap_done <= ap_const_logic_0;
        end if; 
    end process;

    ap_enable_pp0 <= (ap_idle_pp0 xor ap_const_logic_1);
    ap_enable_reg_pp0_iter0 <= ap_start;

    ap_idle_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, ap_idle_pp0)
    begin
        if (((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_idle_pp0 = ap_const_logic_1))) then 
            ap_idle <= ap_const_logic_1;
        else 
            ap_idle <= ap_const_logic_0;
        end if; 
    end process;


    ap_idle_pp0_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_enable_reg_pp0_iter2, ap_enable_reg_pp0_iter3, ap_enable_reg_pp0_iter4, ap_enable_reg_pp0_iter5, ap_enable_reg_pp0_iter6, ap_enable_reg_pp0_iter7, ap_enable_reg_pp0_iter8, ap_enable_reg_pp0_iter9, ap_enable_reg_pp0_iter10, ap_enable_reg_pp0_iter11, ap_enable_reg_pp0_iter12, ap_enable_reg_pp0_iter13, ap_enable_reg_pp0_iter14, ap_enable_reg_pp0_iter15, ap_enable_reg_pp0_iter16, ap_enable_reg_pp0_iter17, ap_enable_reg_pp0_iter18, ap_enable_reg_pp0_iter19, ap_enable_reg_pp0_iter20, ap_enable_reg_pp0_iter21, ap_enable_reg_pp0_iter22, ap_enable_reg_pp0_iter23, ap_enable_reg_pp0_iter24, ap_enable_reg_pp0_iter25, ap_enable_reg_pp0_iter26, ap_enable_reg_pp0_iter27, ap_enable_reg_pp0_iter28, ap_enable_reg_pp0_iter29, ap_enable_reg_pp0_iter30, ap_enable_reg_pp0_iter31, ap_enable_reg_pp0_iter32, ap_enable_reg_pp0_iter33, ap_enable_reg_pp0_iter34, ap_enable_reg_pp0_iter35, ap_enable_reg_pp0_iter36, ap_enable_reg_pp0_iter37, ap_enable_reg_pp0_iter38)
    begin
        if (((ap_enable_reg_pp0_iter26 = ap_const_logic_0) and (ap_enable_reg_pp0_iter25 = ap_const_logic_0) and (ap_enable_reg_pp0_iter24 = ap_const_logic_0) and (ap_enable_reg_pp0_iter23 = ap_const_logic_0) and (ap_enable_reg_pp0_iter22 = ap_const_logic_0) and (ap_enable_reg_pp0_iter21 = ap_const_logic_0) and (ap_enable_reg_pp0_iter20 = ap_const_logic_0) and (ap_enable_reg_pp0_iter19 = ap_const_logic_0) and (ap_enable_reg_pp0_iter18 = ap_const_logic_0) and (ap_enable_reg_pp0_iter17 = ap_const_logic_0) and (ap_enable_reg_pp0_iter16 = ap_const_logic_0) and (ap_enable_reg_pp0_iter15 = ap_const_logic_0) and (ap_enable_reg_pp0_iter14 = ap_const_logic_0) and (ap_enable_reg_pp0_iter13 = ap_const_logic_0) and (ap_enable_reg_pp0_iter12 = ap_const_logic_0) and (ap_enable_reg_pp0_iter11 = ap_const_logic_0) and (ap_enable_reg_pp0_iter10 = ap_const_logic_0) and (ap_enable_reg_pp0_iter9 = ap_const_logic_0) and (ap_enable_reg_pp0_iter8 = ap_const_logic_0) and (ap_enable_reg_pp0_iter7 = ap_const_logic_0) and (ap_enable_reg_pp0_iter6 = ap_const_logic_0) and (ap_enable_reg_pp0_iter5 = ap_const_logic_0) and (ap_enable_reg_pp0_iter4 = ap_const_logic_0) and (ap_enable_reg_pp0_iter3 = ap_const_logic_0) and (ap_enable_reg_pp0_iter2 = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0) and (ap_enable_reg_pp0_iter38 = ap_const_logic_0) and (ap_enable_reg_pp0_iter37 = ap_const_logic_0) and (ap_enable_reg_pp0_iter36 = ap_const_logic_0) and (ap_enable_reg_pp0_iter35 = ap_const_logic_0) and (ap_enable_reg_pp0_iter34 = ap_const_logic_0) and (ap_enable_reg_pp0_iter33 = ap_const_logic_0) and (ap_enable_reg_pp0_iter32 = ap_const_logic_0) and (ap_enable_reg_pp0_iter31 = ap_const_logic_0) and (ap_enable_reg_pp0_iter30 = ap_const_logic_0) and (ap_enable_reg_pp0_iter29 = ap_const_logic_0) and (ap_enable_reg_pp0_iter28 = ap_const_logic_0) and (ap_enable_reg_pp0_iter27 = ap_const_logic_0))) then 
            ap_idle_pp0 <= ap_const_logic_1;
        else 
            ap_idle_pp0 <= ap_const_logic_0;
        end if; 
    end process;


    ap_idle_pp0_0to37_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_enable_reg_pp0_iter2, ap_enable_reg_pp0_iter3, ap_enable_reg_pp0_iter4, ap_enable_reg_pp0_iter5, ap_enable_reg_pp0_iter6, ap_enable_reg_pp0_iter7, ap_enable_reg_pp0_iter8, ap_enable_reg_pp0_iter9, ap_enable_reg_pp0_iter10, ap_enable_reg_pp0_iter11, ap_enable_reg_pp0_iter12, ap_enable_reg_pp0_iter13, ap_enable_reg_pp0_iter14, ap_enable_reg_pp0_iter15, ap_enable_reg_pp0_iter16, ap_enable_reg_pp0_iter17, ap_enable_reg_pp0_iter18, ap_enable_reg_pp0_iter19, ap_enable_reg_pp0_iter20, ap_enable_reg_pp0_iter21, ap_enable_reg_pp0_iter22, ap_enable_reg_pp0_iter23, ap_enable_reg_pp0_iter24, ap_enable_reg_pp0_iter25, ap_enable_reg_pp0_iter26, ap_enable_reg_pp0_iter27, ap_enable_reg_pp0_iter28, ap_enable_reg_pp0_iter29, ap_enable_reg_pp0_iter30, ap_enable_reg_pp0_iter31, ap_enable_reg_pp0_iter32, ap_enable_reg_pp0_iter33, ap_enable_reg_pp0_iter34, ap_enable_reg_pp0_iter35, ap_enable_reg_pp0_iter36, ap_enable_reg_pp0_iter37)
    begin
        if (((ap_enable_reg_pp0_iter26 = ap_const_logic_0) and (ap_enable_reg_pp0_iter25 = ap_const_logic_0) and (ap_enable_reg_pp0_iter24 = ap_const_logic_0) and (ap_enable_reg_pp0_iter23 = ap_const_logic_0) and (ap_enable_reg_pp0_iter22 = ap_const_logic_0) and (ap_enable_reg_pp0_iter21 = ap_const_logic_0) and (ap_enable_reg_pp0_iter20 = ap_const_logic_0) and (ap_enable_reg_pp0_iter19 = ap_const_logic_0) and (ap_enable_reg_pp0_iter18 = ap_const_logic_0) and (ap_enable_reg_pp0_iter17 = ap_const_logic_0) and (ap_enable_reg_pp0_iter16 = ap_const_logic_0) and (ap_enable_reg_pp0_iter15 = ap_const_logic_0) and (ap_enable_reg_pp0_iter14 = ap_const_logic_0) and (ap_enable_reg_pp0_iter13 = ap_const_logic_0) and (ap_enable_reg_pp0_iter12 = ap_const_logic_0) and (ap_enable_reg_pp0_iter11 = ap_const_logic_0) and (ap_enable_reg_pp0_iter10 = ap_const_logic_0) and (ap_enable_reg_pp0_iter9 = ap_const_logic_0) and (ap_enable_reg_pp0_iter8 = ap_const_logic_0) and (ap_enable_reg_pp0_iter7 = ap_const_logic_0) and (ap_enable_reg_pp0_iter6 = ap_const_logic_0) and (ap_enable_reg_pp0_iter5 = ap_const_logic_0) and (ap_enable_reg_pp0_iter4 = ap_const_logic_0) and (ap_enable_reg_pp0_iter3 = ap_const_logic_0) and (ap_enable_reg_pp0_iter2 = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0) and (ap_enable_reg_pp0_iter37 = ap_const_logic_0) and (ap_enable_reg_pp0_iter36 = ap_const_logic_0) and (ap_enable_reg_pp0_iter35 = ap_const_logic_0) and (ap_enable_reg_pp0_iter34 = ap_const_logic_0) and (ap_enable_reg_pp0_iter33 = ap_const_logic_0) and (ap_enable_reg_pp0_iter32 = ap_const_logic_0) and (ap_enable_reg_pp0_iter31 = ap_const_logic_0) and (ap_enable_reg_pp0_iter30 = ap_const_logic_0) and (ap_enable_reg_pp0_iter29 = ap_const_logic_0) and (ap_enable_reg_pp0_iter28 = ap_const_logic_0) and (ap_enable_reg_pp0_iter27 = ap_const_logic_0))) then 
            ap_idle_pp0_0to37 <= ap_const_logic_1;
        else 
            ap_idle_pp0_0to37 <= ap_const_logic_0;
        end if; 
    end process;


    ap_ready_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001)
    begin
        if (((ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            ap_ready <= ap_const_logic_1;
        else 
            ap_ready <= ap_const_logic_0;
        end if; 
    end process;


    ap_reset_idle_pp0_assign_proc : process(ap_start, ap_idle_pp0_0to37)
    begin
        if (((ap_start = ap_const_logic_0) and (ap_idle_pp0_0to37 = ap_const_logic_1))) then 
            ap_reset_idle_pp0 <= ap_const_logic_1;
        else 
            ap_reset_idle_pp0 <= ap_const_logic_0;
        end if; 
    end process;

    const_size_in_1 <= ap_const_lv16_10;

    const_size_in_1_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter38, ap_block_pp0_stage0_11001)
    begin
        if (((ap_enable_reg_pp0_iter38 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            const_size_in_1_ap_vld <= ap_const_logic_1;
        else 
            const_size_in_1_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    const_size_out_1 <= ap_const_lv16_5;

    const_size_out_1_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter38, ap_block_pp0_stage0_11001)
    begin
        if (((ap_enable_reg_pp0_iter38 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            const_size_out_1_ap_vld <= ap_const_logic_1;
        else 
            const_size_out_1_ap_vld <= ap_const_logic_0;
        end if; 
    end process;


    fc1_input_V_ap_vld_in_sig_assign_proc : process(fc1_input_V_ap_vld, fc1_input_V_ap_vld_preg)
    begin
        if ((fc1_input_V_ap_vld = ap_const_logic_1)) then 
            fc1_input_V_ap_vld_in_sig <= fc1_input_V_ap_vld;
        else 
            fc1_input_V_ap_vld_in_sig <= fc1_input_V_ap_vld_preg;
        end if; 
    end process;


    fc1_input_V_blk_n_assign_proc : process(ap_start, ap_CS_fsm_pp0_stage0, fc1_input_V_ap_vld, ap_block_pp0_stage0)
    begin
        if (((ap_start = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0) and (ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            fc1_input_V_blk_n <= fc1_input_V_ap_vld;
        else 
            fc1_input_V_blk_n <= ap_const_logic_1;
        end if; 
    end process;


    fc1_input_V_in_sig_assign_proc : process(fc1_input_V_ap_vld, fc1_input_V, fc1_input_V_preg)
    begin
        if ((fc1_input_V_ap_vld = ap_const_logic_1)) then 
            fc1_input_V_in_sig <= fc1_input_V;
        else 
            fc1_input_V_in_sig <= fc1_input_V_preg;
        end if; 
    end process;


    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp177)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp177))) then 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_123_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp41)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp41))) then 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_191_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp250)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp250) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_197_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp322)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp322) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_ce <= ap_const_logic_1;
        else 
            grp_dense_latency_ap_fixed_ap_fixed_config11_0_0_0_0_0_0_fu_233_ap_ce <= ap_const_logic_0;
        end if; 
    end process;


    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_ce_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0_11001_ignoreCallOp334)
    begin
        if (((ap_const_boolean_0 = ap_block_pp0_stage0_11001_ignoreCallOp334) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0))) then 
            grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_ce <= ap_const_logic_1;
        else 
            grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_ce <= ap_const_logic_0;
        end if; 
    end process;

    grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_start_reg;
    layer13_out_0_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_0;

    layer13_out_0_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter38, ap_block_pp0_stage0_11001)
    begin
        if (((ap_enable_reg_pp0_iter38 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            layer13_out_0_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_0_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer13_out_1_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_1;

    layer13_out_1_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter38, ap_block_pp0_stage0_11001)
    begin
        if (((ap_enable_reg_pp0_iter38 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            layer13_out_1_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_1_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer13_out_2_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_2;

    layer13_out_2_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter38, ap_block_pp0_stage0_11001)
    begin
        if (((ap_enable_reg_pp0_iter38 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            layer13_out_2_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_2_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer13_out_3_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_3;

    layer13_out_3_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter38, ap_block_pp0_stage0_11001)
    begin
        if (((ap_enable_reg_pp0_iter38 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            layer13_out_3_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_3_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

    layer13_out_4_V <= grp_softmax_latency_ap_fixed_ap_fixed_softmax_config13_s_fu_409_ap_return_4;

    layer13_out_4_V_ap_vld_assign_proc : process(ap_enable_reg_pp0_iter38, ap_block_pp0_stage0_11001)
    begin
        if (((ap_enable_reg_pp0_iter38 = ap_const_logic_1) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then 
            layer13_out_4_V_ap_vld <= ap_const_logic_1;
        else 
            layer13_out_4_V_ap_vld <= ap_const_logic_0;
        end if; 
    end process;

end behav;
Zl9CAA5Y1dFl+k+5on1SRcFZumXYSFB+/kdYW0+j8xPwxvrOokj5A91DEXckdmopGqE3+CGZthfB
IvkSTa3cIBBysCJF/3/x/CewWMzd1V9I5tPVRzEO21kNUrk4MDZF8p/QZ4PJtP4YDcy4WjInwcRs
J0jdItpjDbFO7BwjS4e7eYneiXrg4KevkzLWOuw9GgXxLo2Cy2Tj5XZ8mPXu1Sb92paCRXh8DBhB
jNqUSkgVAQIR5s62Qd5Zbc1rQz7qfNsCPRPda58NMuxa+ZXo2yygReAIp+4mrOoCkeV13+eoMf5M
kZwLRPol7Gphct8kk9A+W8G2KNlotzYBu1xDh1uqp4pUU6n2sSE7Kcmbk1tewCGwNrs2BPXbpHIg
FkAbk4ILTPElUDFL9divYS81I5bflEoX/PORW0u6lpMstMy0Zbg0sB60XqCtVNnArUNABw6BvsFI
oevFGjS/CBPB3HipA9TsxqEhAiSv/dAoE8lhxlHuiuTnSxibilLR4fJCpvf1wJyBwrsBs/idWPOK
NLWWH1fF5Z5QfbdSsaem7m70KtrugqbWbJ+XD7Ts0HA/NDompupWTl0UGL6HXdrq5jxyQ9waR03u
R3WHHXGkk8wfjS8P1usfhwo3mwGieCdF1QKhPpQqUGp6SMruPG9TOEcDGMWfmouZpq2kyPy0bPP8
THAeGkCtY3CWuVXlm8yMgmm/LnVtPIrRXrsQHPCz1F+vpNwOf9/rdsOaxXEAknNooayG36WmW8k7
i3mxYZguhORxmPXJXgqbePHKnWZ76xHbxU9df2wE6RartY2nasIG/EKEB2AiQBH27M+jooSCeoon
KY85AIXrbUpuNGRXy8FXjG7CwgFu26dhufPYCBZ1ONqMJQDDR9PTMY6szeazolNpftJPPKyO7iLq
+avX8haz7rSUxBvAmxy2nePj5awHE99gF4oMqcX3elz3PURf5ilHvueRNx/vg7CgTMu+k/L7oLm6
JchY4IdUmKpiT1j46Ydo9NCSDc2Kd4u/HwDpEFLqDbNmfHYSa6z537pGThOL+2kCzHz2XAOD0TUG
CVUm1a1qLF6Xcw+Z+RFXzsiOsd8YEYe6m3sP5Vwi8VV6qQJOTPIW0kTi0ybAjaTZfpdsS05qhwg3
U+dNQBPwOwLJGkSRIx9/tpp5AxjyAKB1eYpsqGTnlGFlc1h9vrJeiCNQnsPj5mmJfG4XVWn4oldv
r3Ljk8Ru8bgi6a4u4JhNNYTbqLhPmQY3IMVqC9DR7RqGsFZlRaCBTAdMCYZHbNPPnXo67OtVPQk6
6JUKDA6sPA5cf7DeB25grNd8BwiGhL56st5UXbHEA5rTSVuEXy2t0d4N4Gvj1jgwVIqy2x0nKJQo
OEVtVybC7v3gZUdPRwnVr4AZh/U0wspJdlwHVsXBzqrltjZZSPkijhOtZbRF5MrOoi0b67aUQG1H
2g7gou7yozfyqXKdOh2c+5F3osYIoaEEHgNaUZeIPG+vRJ5cVJ+LC7eND7PWdBdRIsbqmpCz5xrD
8q7NzX0640SxZZBPOoI7UfCkSui/rf+4WYbuQDDQhcGFp6rRTz6jL8hKySevSpZ1UG52TzkRNyt/
89A4LHmIuiJOqK576qpSFGf3IcLNc5To1W8nBT2VitUeSgZIcpBGaX8K1ekBQxnB9gBbZzjHp2uF
TBdl9K5nfcstNNEPTEISxiBZk7wWqhWhDQZfxgC/IHFH5OTxViu1ngoU2PVYWIUrLv75YzKvJy/g
xTrCLBZzuw+ZM+ConOAhUdVa+RfE1un4iOYgpXx+JRkCIxdgDm4k7mpKyVNpAvYeOf1wFZBSlpA6
GTHOPU+YuWrwBYI6vq6kbIYkrQuEa5w+QjLuFFHfTcm8nBheKOSZzbH7Cq3Kvzz+J0mJJVwmsk1T
fV+GnmuvCNV7r43vIdC849044+mkGb2ik9M9eWlldfYJ/8OBifDLaQTZQ6k33+gK+8b+c5p0JLAb
O+NCt1li4RpobdhT0eFWo5xXAphZxW3EXMRs16VNB1UEX6Yzw6CRwnmyLuKuTgZdHSSnXeGw9VIW
9L4PGYJxXBq4NnKoPSNFXQ+aJCk7N8p2TUCx8KnMFWTpnGpjoOzTcBGU2qst8X/FIwbSaEqtGH0d
Ju6+AbLziGHUv1JGXmbBT8tlpUoKAmK/Kz/LuUiYvguLEoMS9DGXTNt+nrruxNh9h2DZ37HVTQ9c
1xUyNDwO0MUFbm90kGkReEPJGahyPspLdpqBf2HV7NwrBTBnBz0+Cj7sFGHiLRo8E1ujqbPeFAp4
y3fawVAYrDZip8LcV7UcRE3D7pPdQ1KrfiDciXW4g1WLR7M6s+2lQMDzTraCVOAwmZMCu7ZkpTQU
2TyBH2XYyePdffNmZ9mctK4RPKxGkTuTttZG4VPb16avBph/u9Py2jPc4A0tJ17UzJgtKXkOecIM
Q8AwGs16OLFBKwrxelyZXJmA7mEAWfB+yNmQhnSOT0Ktf/xrFTJEVYNUOXPYDZ++Cq3TIb91KG9V
CzGc3Ez9Q6GQn4kCT68aQ3fR8bPa1xF3ZO6azXc6cmUq+FMBIIkAdnGVllIqNTCD3D+Vk6gThwt/
QR9OEvnHPpne7AJWHjTB9QVdopCsbhVgiEDPvE3LkPSadHW9IBDCCp0YpjgE0J9gw6r1w+2NKEwM
/AdyxXQedtShuWRBbf9/1ejAMXqD/RttI1u5PoaBKNg40YqmNOragNxDVHb2FZut4nGMSc0BTvwe
M84tPazeFzC5DEuCuxM5bAmXt1MjNMsDpwECJGpJ6o3UJ8nPC7a0MGif0ct5ulmCv7LFUH+xqQcr
6BoN5l0Ol0bM+kYP3BfJyNMl2gFb0Z5QG5Kky9RtjpG+cn0/yhqNW4e3PW1v6/OWgVGICfXSX2hM
cAF018CqnaZ4ABzBjyqDq+XpbK7omwerXutmsCV+m/tRSJqx3WL6GnM814PVNCuUDXGU9TpAyOZ6
ceBBRcSSPSz/xv5EWjfWkUlHU/2EUBkwpMB/SMbkfmjrXbQlpFhvZK7a9Aq1vEdB3vCdm6yN6N2h
Utwhk4d/Gm0NRJHBdUX6BWICfzWFPC8gVL8uomLsXujnb+UavHCYQlFOMrsCGlUpvpgjWLqT2Avi
A97GvliqK330304SuE3d7fBefJoThJBKTW0iTMzx2rSlT9ITnkeQk4C9Mr4e+5UIEbt9PDAHeG2C
72EovBfF87aijuGUS7fE6NZy+MdAziZC/nEbhp0MB7YEmGi8dgxcn739DEx9MjCwn8TILTtK1aWE
pfqVILzFEed0yb/0CHqWAhdHzBS66XoSYZj9pNlDzaQm+NFRR1FiatCO0cpGL+L2hQS6YvOmFMdA
LpCsvc0tmVTiPkPNrkeKX+5GGEjgiAo63AsGMsVd2CidjfrTxlC8FcceVjhwc3PRmsqq5yCddCpt
R9obpMc6WSidCWHbCOsXalFfzGyLvG9aV9/UptpiedJIv0jvVW2otNXpCd3GbfC+CWugG1FH7QFj
pQ8B8K+i9MQLBCSjlgev9m+/osxUNMSbdOe5TUhvxrZdZyVaCMfyya3obRvHHno+GmnP9fsC/9v0
Z5E2DwEN0ehx+p6zqTqrxdEZ6P5g5qoDoPZaMmsJfr779WeLGJ5pvqPIxPeXKof75cf7R2GHsdSM
la9vXSoFG7KH3HMX4acoqBnK+UXvLCs0qmLNX3OwGfMB2SgXqN6PA8L888iZn62L29L44BjAg3cL
wP8qTGu6qIC7tlveloyKT9CUx1Ux/EIlQWry7e9SAEhHBJ8NlAlZPjVclXqRG/KZUYZssxF1TyaL
CsGt5nm3Kjy9/AIw6jzPLnuqKrT1qnCR+oqFw5dgplhVPnBUwU48ZYJv8PUb6zW3xp56qyCvdQTp
su3R79oGf2uR6QLR4UKk72zBODnWljKd+SDqhfQIARiVtYtWpJrlhoPkMu125wJ66re/hTByrfIX
aBYjXsi6eTjWoPm9D7pZkcY9P0O91266P6P/JwJNsQpZJURmFiTFnkzR7x8d29pGsQmrLWCeu31D
NOibZRhHzN7ahm69tcN2AZlsGHC4ed0sJcJjP9NogyjXmZKxhJfkpSgvODGIbL2hbWkC/K9oCrfi
TNbW3VwNBZGVWZriIPk78deHD0jg9YlgbhZ9TYIRTjb5QelhVugvfEr++JPqnYlizXYFwRn+K+A7
hTG+3/lEQsnq6BXtWWlbMVKkdwWIZKLHN9Mw61JEtdcq9ltF7+D9aALgQLHWul3TpZrueV1QmetW
OrujCFFFJ9ofDGB6uAL/mzfCaxaHH93UakvyRHPA48yHdjDeoVr+cUHRSyb7beigCqhY82PiU4Mw
ZCD0R5vIOIi1goNN3+ZoQAB5tmilBozd7aTe8B/JfonBc6BoIQOpPp7awHaeuvpZEWMR12UgwQ14
STfIY6y/bSDD1m+0Jx20q0vN5KnYk5dLM70j0stfPvp9nDtwlm2NlHw0oVSlF1Cb+UZAz9+Nct4v
WAxDc2I34cbPhnXGuKLCqL5tdwrMBHgIdZBvWZ2swkytAlX+yNH8TJ+5kitsk8W++434aENPFnFb
1K4JbKNYnVOZakrf5IwCnojF8ydQXrULiaZo0bKWb8AxV8kZzGqmzC3oRDXxI4ATv7/b67r4pvr5
8ZfJztgexQN7cm4ZGJPIUO5FZuMOjj1nEGhS0ywcYrkLmZO14M5WLJR7FLc4UpQOTBImsIvIxLf2
XKus7w/pFJ0jCdLS3Gc+JRlGOQLsH3KG3AeC7TMJuVQWGm08OvqqGPoKyXM5VaGVBeHAYjb14qgL
KQj7g0t5K4ZEREGS7t7uXJyfMVejhBZnx8F26d1qnYAT1k1iUPd5ES2jrnT8cMobbOFwYYcOBg/1
GqevWc1crCKZvfI+98szQE8S2FSXfWsy8r0+DVAc1tRqWEkfn5zk8fbxb7/cJl4Z1gyAeybN91Ai
D/la8qcDL2zPj98+pIsFxlie8jEaLjUrPRIP/BGw2pGGJZzXrv1KDBbjyhfXaPlZ9R8j4FBXYLPs
v5ra12oM7Po75wRQaadjQg4mEQ7jNvCVJg4DLwDMLgdvTQ922xyxf/PUwKBZCSj7sxMH5L8/Iwu0
M4CDJQznzLQKXAzugz8n/WxfKHXqfkeHuYtMhbR7BCLSnmC3ai9nEqA3AN/kADH6RDKP0meBvG9o
oAJ3CwchdzmqUbpq85WUYm14+vEUraHgh28NL2dxzTOmTgxs9ODhn+m+vHdEH4E6LhDJbuarp4uE
4zmIu9ChSiWctqZk3gmOOuHLiZ5CxaxqBuMhEh1kY0Grt6ZLVDDBRyPxMP6ndbfrMZxnyC2dwcVy
snJjdFWBDiJw8jYNAmtCkRjdqcj8Imk6nWqEqyPMgedUKWQDIQRbWD9AIdUMzAgUp90eIjOnfmWL
mj46bAGg3+Xwa9gIzJwfSSTANL2L3GiLegKLAaGmz6fboKtEXrVGaz+1K99wm1Ha62KsAukbKUY5
//p3e+ZJ9rc4ykB71dhKQI81jcxYh9X71FJTqqho5FEp78oAigH2A3jtYjxsVmWl16Q850PgLR0C
xDgLuzMIc8idP2yS5m0bWAi8KfJbRLygdibI3uvE8aHJF6IaFMw97bJakQcSP9pVXAerttPBCKjt
meJq30eFfV6AH8Tzxy8RjNH9Lf01dP0IVzsOx0l45KT8Sgy7Pt9YVoAOlwO7mqaMsxQkwEApBFWG
si5dqsy6PCUKiCL43N7RCdmEMQ5WaIyG55xYWCnus/RsSlNDQy0i9hbSawr13CXiMIJ70sf59INC
ckowDSwyt1+Qd87x6z4SIY0KRg8nYryIyLcnnON93Dww5Oit5YB6ziebtfgRkLcIzzoCW0MSJioz
6wNbouxPN6+DQWoZ5GXAmNXL36xupS+xAu4eoBmNTA8ZhowXaKh0kClcsJcLL6kBvVizKPL+yq04
DwfEJ0103MhhNvc1fCgeTF05mXFY5Mi5/biXw0QY1yeKN4mjqED6+gbiseMCLCMn8thk5bNDTilu
wEJXV/+ZfWZzM4fyILdjLkGgH2cW8Pq5TvYTwCBeQ6kA4/E/ZLINJVoxuwwfNcPq5WSGCEObm/Kr
k4/ETrQjh5M7mvZn2kGrF4IgSS3riLHn/0XRSdIB6lmE7YYldRmuXG1cPZY1dyUa0EoVB/21iYl3
efQ4lLNZo3QCKf4JVB2unW0IlBq5MQ9u0NRtaGTpXDg9lizJohmgSkrfArXu5Bc7NqVsTOJ91ao8
JRitM8gLgUrtmps0q3uP+A6NNHYbflfosKkTT7CHZ0sJuHQVYxMC8mNIX4TtcyJ9nXjIj66ZP4E0
+rL8mvtRKvf8SC4rXAekXgo3mEpWIBA+dsT3RYE1GO7Jr7zDMLa6psu6uPTB74a6FrPgNh9j3GH+
V8HEesYbiI/GZEk7rwXWbvPF3m1LVpiu+ifXp7Im5oCSLYzp4my9BGvpzPSnth+sRTrmHKBr9ncy
zm5m47tVxm9mmfsuzSAAZZA/PoaaIIJiWs2nEwBwOto0SVFue4w0VDeiFPl3Qzz+R3VuMwgK6+Mf
zxBVZaNwEHr/MC2m97+/jJEWJ2TeDC90i6H8zvaM5Zvx0s31y2hHxyp+SGeuRsEmMQymPQ0WXU08
5A7TDK6xPw1lxZzR1ydJvZCVH3UY1bME3HHqy2p/WVfnmhGTdk5OJotaC0hCVRQt4lVxtlGeElVN
TNd95TBUZ2S35o1Nt1wDDgawyUcjba+ltzA0dXzku+grfgpJn97JU+QDoDzx13zETtHesmgX8iEd
iQ2DtabZUEVDA69eHZEPJOyH0w8xXxrxHYuXdUOfrDTlMYb/mBqnyTw7cnLxeyDM0pqY8V/fXAXl
x4d4xsKrKz2W7O11zBfcY09VD9Zp3k0wdhHhmqikqO8HQXmcF+sWwmhLklxfA3VVfFwVO9DbBjIH
pvbEdPJ2Rej+kIN6yJgwFnnMhvoAhd+WApTXQeOBagxpZxjMh9FQy4kXY+h5etZr9nO7oHlcr8h6
pIu31D1L8BGLTopqerTwRUEwzcHWncMbMjbsPZ4+ljYJZwvTMB3csnP5xvrGHLYgSGgDGbYIwSxm
Ltrr6RLJYd/LKsRuNT79WCQ4X8BKAOfmxn80Q1eXLSmo7Ek/R8B22gOBbepNE3uRZhoZL1OgqW6b
/v0+nYxtG0FuWdZX3q2mLyWdtLtDoPv5hVRCody89vCRCyIkocXtVOlBpBIJX+L3L/binTIp5WTm
YXGiWkcoWrX6bAK2b+EjtmLEZjihd5bZoMf9ZVpkuI/5ramnB8OSijrGAYC6WUSObOb3RElyHxo5
J3tix9DO/kGy9W1fFCZeb5P93ZMjSRk4EFCSrmKxc1QQEIFTA2lonIuSbMsuryZRFpxdh4Ropcuj
f4QdB1s432DEnAQAL7EwDUo6q964osdtpgQmDxef9Fyl/kp9IY/jagwGr5VLBSIQHJTJJzvepjeR
I2ORFtaS/aOB88xukwb+DW/lIP5kTjla7S3tkHb1niye/nDAJSAi93okEz3K141UOE+d3TIsqPMT
8URal3gNs3EC1Ssf+Ezv1VBIY05NehEGEB+/eA9CDvvFQtNrF7P/sy+0G991aZzYCmYOamt8Y/w8
TnPBWHu/iWEko8w0HWXfdiDdsy0FOmHy/MRSBBO7M0y/9LhEoDJtWn1ftN/rr3DyjiO2tYLINbiM
Pe4WghKl/wdDh4bZZOtXWGz4bKV777rBk04AfpwdvlYhCFNx9GwzkXi1NdbLcFd97Wmv829+sB8X
EiIYn/8l3oaaUDK4HZQPHTl+LWnyeg2ahE130DucxxBHN/uEKFZ66KBJBU8QiWV+mIvPuBKsHdpy
5iYs7B6e+gQWQ9rT/6Z3Jrzs1Un5eDDKylFqF+H2OjGlBqKuTXkcIteuDnHDHz6np45NOMm1XwCs
mlqdO09ems8CIOhZkscPWC+WkR/OeGLFsEaUX31uh0pspYrh9oI6gzWv89FzWREz4vW3zpKo5a/g
YWsdTCpaXtUnOEjVJDzd1z+3TtVYQCRr7gsyt0opRwEBhYUKN8/J38WlasxFAVtuwoQrAiBSdcTa
YMUWaP+ZYY1tzeGdT4ue69Y+jhdoYEBe9PqXWIE0Y42K9Yo5etUWmjxTG4znkj8OTRvMgTKUdRMu
eheNfjhDNn5MhiIdLkBcOj6NK7qlItO/xQRBq3B33PFtptfjb4UMpO5DaOnHdbT9MJlZzMvD6ZR7
eKrsO9sBgRVAJivdoi4apB641bWoRIUtEELIOyTL5qfVQ3rTCFPGPsL6QZ9E7QInUHFF7JXYQhCx
SRFZbCiXQmQrJLpNmZL71TXc2OpMcN9OU0Pm721hSO9ZXRN4O1P6Yr6vvfVmPv8JntuZIAprtglA
U0A8xRkhu+0MkW1xHK8If4mPLUz+hpBaqsob3Fh4/ghfxun1C8MTgdwj0o4dNjpilx6W33IlP2kh
pPADm6y8Y93uwZKBBX9Yji+nihUQbRIl3nH3H5GdIbbG+niRdgn3lQsaCRyWbyKIppIvsahPMjLD
kSDXPHVA1kyAh5rdKPfeBL2SDnlX4K8oVYplWKkcEp2X/syieN3NmixLtu20NxDNsgQd59zZ5KGc
K+pAuHGYwuDYeNpJKZIQXkyyeC815BYSBbE0l7VCodbSWkPToaMH+2ll8ninnx5S7w54Ppeo8M5w
Z1VgLaLgSucIH4kVnJEUWH7IO74E7jWsxUwfArFvgUosfyp1+PUy0U5jPeu+vr/X9W6BNFqAS/mx
yRSEMCZU/KgBnpVkNJuC84PoLfsZfeeO9PgDFvWeJ1hvd4Cro0LqAa7RCapMe8+WLi2t/y/8lVsL
5JTkRdPpuAeGYChJQ1NFZPpJ2YY4TN39QO2SLM7z8cmE0eGnXx7SlQObijI8LXWLz2jzmHT4BbTX
pdN70HtxGI2+sE8QQ8efHBCpcSKoOexrnqkpcrniVhFOuMQKlgTId0l9tCWrDVi1MvuBITdx2LPC
uln/VHCktmkqVGb+j/GkfCogaG3d7Lc6usqsQHT5RC3zKxkbj6S0RWxCAdzQokNVdmg07nZaKDoc
3JpVioTlHKq3Ihm5JbXaUjjn2iHMd98ZfbMaObk2i6ys3Kwk45Ro9ClEi7qFzoOSFNiyFAz03I68
j04QH0ksLw1IlCBC9ut/s9o20pzgTTXH0dqCKwzo1O7Kw5vL1kw0+5cf++XFo+K/ncY7fOuo2Kln
pVKtwnTxYm2QZ0wUTow5yJZlXg55xOWLMZoOprO0R49jApN4j8GAcje7KFx+huqTINcQqd2+Vpst
qCLTOGBoeQvPJN6o4jpJKoPI20H92woCoC0gKwaj/kQ04XVmOT9P+sVmCcZVR4wSuES+q51zfRF1
TI0gQ45WnLxG2AnvsibGgYlzWMx8NWV/yNuOxBQaGAugCnyStE0fHJvVTeRQ0P44wpah2sHuh075
H6bJXFqalHhkxsatjSTsyHrFOZRwoyvWqhzuOiEiLOrehKrK4Z32SKFsbUOfbgxy44wiSEg8OLgY
joac2wnF/wkuSAhbCZf3afCpLa0NDbaZTJTsEPZXbbpjzZAIBnx92GUkRtAgtgl6hWCfdtkcCCDX
ooSO5EsHdCYtabxFNc+DtcZ/IokqvitFh7IuQOPxF/dXubYLgQzIrJGZz/qrClU4vmvsV8H7HRRh
/sfLyNACrFCkynfGlykVE+klpuG2Pm/1dUIgbvr8TCUPaKkSC6Vq21XkdR37GoMKWKcXdLJW5qK5
u8Uu2iu2eoYJehXilzTNmtoPTIwc2SNi2oWBl+jnIA1fsGotVpW7LUu2x0wIHEmdYVZ9214oiVl0
Dvs78cNVnMe5i5cKkylByF0FpQBgGE3gTkOfYhscwk2LmFog26BoL4EbyHFK+BSGWFGQt7+o1fpN
LsiTfHPBcgBmV5CVTFkopM8F8hz9ThyYnCnO8e4mxO85C9PMeLcZ1ke3/jaOCoawQXEBEyXcyjbY
+qMr0ivTZo3cB/TKc9Cl177hKYKSupOxIoFTDwzGkJ79Ce92q8QnmC+gcYo9ZuItK8u75ymDGlCJ
Gg/qf6Y3ordB4BZBFe7LFn5dFFQaM3GJ/eApGAz9A5Tg2kxRvDQh0erorPBJMKZgU8Np9EK1jTKJ
Gl92fbrpb2UbrXJzWpsvUPPLPUqMg3AbBcP5yh2b1yxXJj8QtsGOIlO3MhyXrLYhp87FdDI1qdH4
OksFKEaNMEYNymmJ8QQiNBVtCWoQoPtq9QgKd6G66p3jxj/wHX6u0cMNzj+QIuG9hWA8R9/QsUTm
2I6jwiW9BjcPlf5+6IoFe8Ph1U54/HdP9E/6yAD+b8gXfdQ4E4V9yxYYQbZuQwCrRdms8qkNTAqt
cTt6IiQdZFe1SzE/w89xWpArDhVG3XdijdGoJTUDyJkzfonPTGvOynMN9wcBxTQoNVGAxDpTPpzU
aiJiNS8rm08HRz+bbaYvg8KY3BhZ6H2dI9fzxtyBPM6DiG6UAvHT3xRXlH5PzsXEGG5M1XPIgj04
SKyxkcExQwimxYuyq1wvZYAy0v+H93TTxTOzJkCXdvxQuTnkIS/fqCkSKn0rMXLy3Vi2V9sbdZ6b
fW6fRGgH+lLHXRVHxquyc9zm7PsorXMW9/dZDeEI6vSc2SEICtpidzkl4iLEG5ig0QL82wBtiMH5
E3qQaKfEB+OHWlkbssKwIRWDCUwuvcRBtPk9GUisgFD8PnKVYC9gKxm/RafZlP0JHAclesiOO3wN
41L8SKZweiBZtb3jtifEor5Nh8blClF9hxnUKVDWv4J3ZD+p3BDAq0/h79rFyAx5vZvQbgy4FN+t
kEqdwBjwpshLElD+HVoXwFLQzIorWXF6rQl5NF5EtMcd1SWKfe577r+5yC5bV9IXPlRllI7ES8Ne
ViHIiNieWSPgdRJTFBFY2i99rzu3WQ6FByk8/Q5fb673whRVCemM2+paQxvJwCbWkfM0Z4Rc05Ow
07xfzNsYxZ8zUcYXyboDZ7c1n8QJeoykJLdTeOhDt8rRjUZJACn0MyQYf4lXcie9g6iKNHfTB+kq
bHcFObk9toOfm30Pdc7fH1XydE4Zr3HbaZpgMZmm+q7mBTtz88+TOiSWWwh/KZkBKWMmw3Fy3Sxl
cPvmMI+G6nclMnC7LQ6iuWGeqCmWqOC4jiPjBk0KY2tAFyCyyFfYCCBt/0A7xXqWga5USwmD6wMi
zErHuXLgZEU8TJAJGeD673yvyhjewiuC3QhZHdz33jHSwRLoofeUYznAOLvjFT5+vi8uZrVQ362E
7zDPQGLPE/4f+9Tj3wgoKsV9QVyWC/BAOw2oGetKvw8sD3lFOC/FSgbJAQ1NUxAPD7uRfOuMA6lV
mZR5I7r98jLacBqj9ySGPGxM93NP4zVoxmJvDPyaLsArin1FdOI6cny4v8VEbH1ksiy/TOGYMOSj
utAdshQbRkzPKPGjMFLbvh2OkhovrbYOeVoylmsclmhbNRDY/U95aus9tBuD4Qt7tLRnUgblXKtS
p8LIN8VNLuBy4TXXgGZRQVIztjoNcjFFf0MbIvfWuyq/9hcrvg0oIg/LhCn6bcp1EiVd1pUH4HYD
DSQjOf5SVEzbziSmgY4B/g1tXQkfsbO9ilff85z0FWaJbaXtnzy2fzO1aDC4H+A9z49OJ/aHHcFm
tPDVaVk7H4H/SKLeXvdwS3c1/L7AvHojZ9TNdQFCIgQFdo3wFbHoGtKWr/PPrrRGAPJ787skLjMV
JLRtkT4IE90SPmIMX+5KrhFqLir2bdOVCejx5InuQyM9I/7UAwH7z4OH6qEo4JLvQz93sk4btWPJ
RX6LZRWVLh+qd3AR58WGyXrghFD65NFCXRwEIr+EPrmzLbc0Qt0EUzGsPU6yMbgWFvtkH2Iz2u2q
9JrbfbZf2q8yjLTRuytrj4euoiEjqGxTU38oGbtsH/CEGOmNhXKvQhVwZIVG8n3ZPEqFBNrsVpyO
KvfPVMDwFfNhynwZdZv61qVjxvdAtx37DKzq8R5hlz8Fl3XVWoMIYOckbyBca9SCGqWdegP8Xv6Y
GadyP5kQedWOh4XJ/vLVHr7mf0XTgPjMA19AnWDrSgFm6KRX/jRV8ftRee1OtynqI2zBlwgQPRPr
24cKmN+cSq0XIj3aGng6IWUb8Cvv6JXMbOl79uy1tyuXwIA34gPiTvBK8nRjfr81UcbLN2NoyOYT
ynvG4q9xycYVj/eUk6wAkT7OHQibY9lAqcbpqIgJsxaZS3MkHh/m8zWqw18YkyvEBzHZ7lTXbFHt
pTMLECBcsVCFvpH+XTHbdrO0rNcQ8foKySeHwBTky5OV1ZfRW+A1spWmLbWSGGYhosiaOI/ATJmI
ZRcMwjjpKnDBsvT08KtcC9W9u8iEW5opW2f+yiXrCMnhUEe/6S7W8E+lKBlaRhs8wxkVsn+VwQpJ
7+toJR2GT9sbT+Ph3Kz3vpk1IhTxyabFiETLsp60eSvYix9DzU8+1IQX2JQ4l1cE2IB+qsuvPef+
wBU12ksXx0RKXoE2EHxomCFDb0KhD7mHapHJot2Llbb3PhsQKdcgy6sZ8ueb1NpDRVtUuNBC5o9T
FUO6j0qQTmBxVV2GsVG5hYfHFYXJFRXnkZwCErPuuZ+bTYmuhVABCHDTakZuaMlFgVTLHx3NLUSb
XfUxd9yHJfiEADrQOLSljY3jgsF6UkMMMKXoGlvaSNvbdOXvQapQ5RWOn4RCGBwjaPg47Vk8BbT7
1lElDyisZCfWVCaxl/BeBBKQVYthtI3VsayJTi/uvUoUdj/jKT1nbuulu45owmA1ZPh4R9bXBsoX
JrSJ6Vo10xHNsL/bolJxyHywU0t5uKc7nTUfa9aRZ1nCrt4/AlsrAWh7jyZvMPYRcadLzAkqa0ov
oU+k+Fjz+rwsM3pTYfLTeCSEU6epBUzdNkW5Pf0erzJtRzNZU2uP3zE3/TYDuc5iENepXUhL/JTb
9TJ8RfdJ2ZdhOFhGIAZPAqU9bed4dNjvNnhT7BNEODq9u3VoDMwws1Q07TSM1GFK7AjHNB9f6jZF
szwiemwlr3BbrnZzgCH4Bxjf11pqdhqit0XXgilEFjTLA3/XtB7HV79SelwGmMmc78O9eMiki/gz
+RPgVlWkUvtXXELUNaDujFzhwzV/TFtEl1qX3EXX4KVYgpMWpust3tBrqt6yiZymPkTMYJ8zn+2p
xGsPcxAb+Wy9acRCCw9SeTX20R01izpH+JOvAocZtuRETb1cILaU3fdLWukrkMdgCumMMD7aSuE1
5QB5z2/2LjfMML1RoyuAIWYjbfui73DMoHPIKzhCFL725dKdF64alieRw5dsIuvQFo1Kv6Htab5m
9KrjH8WsduLSr8AqvPuhuyEkq//Lj6Vj8yv+aTeNPNKH9DaU383ReqSd1gf7zk7tKB45zD2pT2G5
h+rlHTZxCIp7g7/vFkGlk5MLSwotgSmpHKR0ehcwS/I4+BIMt6yFyx9pEqZQLOqFULTtpwoTJRW9
mNlfmHIKpPquer0HL90EdZ6AvsSPioY0RhzBg23R6+570yekysuXNEiR2SEDb0AIujMbi2y9Y42A
IvsPsY/bMFKiv2J4QAv5b3AKkJWnkylk2rHrmGYebk/m+8p2V4BpWXuW0VxFxHPSfWspGk0aArbm
R8PxRTbzC5PN6OKPdRDDlrfe0b3KFGUIh5cDNWtvvv/5nelmGo9SWOxBguI5ILY40PlspyQRpL1c
vDmqF8LJDHR7oUTdMPlphLzPofsi4Ez2Q8qqsfLxfmo917m3IL0a8dBsVRVV5hV2ycgNrnePlV7B
kQTfEcZeLR23bCmf8+WFfVy5Uaej3aGispaRPHiRWu0xYx0bbEt5Bs9+MiqzZLmeS0mdPbiJfdae
+t4Ewp5yAdxXbY68Wjm/gJu0iFe0EMbrcP9snA8PE/HOa95tapx9eHbIvNKX73agX/tniUB6Nl4P
35XHg4FLD+g3iiZqlB8J30jq8X9uj3JknwKUPd5vm2G+glWkLBn2kjVkKWoLK8Bzv25NC5f4HWWM
AlPqyjMqN+NlteGkg9qKZodiiCzirjN1ek0lffIAtPnErIQkQKV9fMXkKCNQNsX1/nGoYib2Eomp
4HiiF1TDTVHvbFxWSxlwJVESf6jMTu+CdeaI0uHz7KvP+n1E9rRfeLBmBiWMaN8NsqWMN8UKPaXT
Mt5oAqcSkHUTsaLqFn/oZTpm+fix2zdPBWy5MhC+89qYo6QWWYyE/J00LM02VMgG3WS+fod7+URs
T96GK38ta+USeIls0abpu3uB3yfNUqOgn0VU00EQdWgNdYl7+cMMUAoFbqZaltGFZ8EpPEHP0C3u
Wpd7NlG0t701HuCc2h73QoX4TdG9mfAfnz3KJYbza71VQmzYGMtaLdnJDWM3IQETh6T7W+PjYXyk
VQIJahXQ2f4yCqhfh1gAg8Z58yr/qMp0UvgsrY1FAp1giMadG5SSmpuBqoh1lZHJsa6KCZYdm2d4
xH6sdxE/Y5oRHnN1OOfD3zRrGw2LlLTiUjmRV5kbx+M6Zfu0j2PjMdgNzg0isnFPP7fCkid0N6SD
Xw5iM1g8JHjFH0dmgVbaYPfptWYS2N988uD33TQE+89yDNIDW+TQJUy1OVh5gJT55uv+qbEdhDGu
BQXTFhvy1mEvOqj2m52LB8GOTxAD7TCmrZzsXgJjaaU1p6/uWSCRy7isGXC00qqSPgizDeQMSOQa
iGp9jyWmo9To8gUCFVPKUg9ZWDRJG/9VDTDZnNjvyp5lMxyQTyYt8pn73Y0WjyycUi5JZRAzQJBG
mcujobjWC/EEfYjDa0bRv3BtqcAUJFSpiVc8uPyveBbi4gTA45VxiRGwcPCPGmL6nvA8Hm842SYO
HZDI8TfyiJ/UlbZTEyqFGAhYt5pVNs7yJKU3Uv1MBknO6Ar32GUrz8um5qmQzCbt49nzAPtTFTfc
lLWm7oAzfk1kxhlanxOl53twUs8XBsnIN8QPWbOilY6PmPm3TOw26eD2fmLMV54n7Or5Dy1L1UzO
1JRbzMr2A20p8l6H49ClIrH4QIY2Clv1cn544LFeyG/t6lHY2Bf1+rTZDyESDLpZSQrm/nTH3Wkj
zVgIiS4rC0WxJ55PzlrEapfO/twD/dnQ92eyNV7vvvATGV16au5Tyl5QqPMY7seGX0uEeCKTspvy
2Sp4BIWgR9f4XVmnTHw4Ysax0Jwv7NRs6BvFNDmTkMItWZHbMrybQOUoOFFHY+GElr+SPBEdsriN
